��   ^��A��*SYST�EM*��V9.1�0214 8/�21/2020 A %  �����(�AMON_�DO_T   �$PORT�_TYPE  �@NUMJ/S�GNL7 L�$MIN_RA�NGI$MAX6rNOo ALxp �V�~ �COUN}TJ��AWE0�8 � $A�W0ENBJ $��G1LY_TI�V$WRN_A;LM�STP�
��E�C�.�W�TC�
J�AFT�_CHGxAVRG_INT��{�SAVE�YP~1ER_REG��T$WA� SIG6� OP��_VOLTS�����AMP�&A�E �#E_VL � &D'>% I*f$� �_ANL�  p 
$US0 S_CMD � �PRIORITY��"UPPER� �$LOW�$�#$�FDBK�"�RA�v �!SQ_AVG��#�#SD_� CEp� � ��$ �� � LIN�!$A�RC_ENABL��!� 0DETEC��!< ELD_SP~�$PD_UNI���!92DIS�"�I�D IM�#���  v1WFt2���CF�" � �$PS_MAN�UF �2O�DEL�5PROC�ESN0�0WFEE�W0ESC�2�2_F�I#1�1�1�7T _A�O�"�2I�6D�7D�C1�6L �"{2 ι CNV� 7 ?  $EQ�z,xODOU��2?@�TBd  �$?C 2 �Y>ADD   �, � MM�!�$D� ��!?2 $F� �B�?@7	JBSEL�10_NOJDAT�A_s@�@ �� � WPpG
{M
�{"�AWP7 �L@�L
 �WI�R_CLP4 �L@ASBU8  �H $4���R�4�YPRE�F� �U;A_ECU��  JB~ �S   $BP�EEPf#}!SCH>7 � �!���`�1e#dPK�*jFREQ.gULSwbSP�0fg2@y�!hyb*g�F�A;AI6 �ZCo VG}�hp dD�e�e�`P�	�a��dBVB�a�ZEROy}uS�LO]R�`NT�!P��cO	U\93�L FO7RMA0NAra�0�J3	� D�c�QWUXWSCCC @P8JU\�uT�IOEX7d� �A�Wfxcc�pS_91INp�� :1�UJ�� FAU�G"t0LO�0I�PD�!_�G]��R��A�p���STIC�@J�R�OBOT�ADY�H�ERRO�SE�d��`S�g�STA3RTE��!TR�0F~��CHDOG_�@�t��0_ACTIVtW��IH�TOR `OCOLL@�ӃC�0�1Q�2H��qE�2� ?Q:2TA�B�0 =�f5)$g1��RE��@92�I� �1R��r�%;E7��S�!S�UC*�N3FAILf��DSt@��LT��sABXP��NRDh2N3Px��RS�0�Y� N3�Q#�+3����)D�)D�)D���S�T�`3�3�3NO� ��B���Y�̤�0���R[2����� 91G�.�*�.��<�^� ;���-���.�S?�0��0PA� h������/HOUR_P��o � ��SE�0 �T<�:1HEpP6��GA�HPZ5�Y7�QLENGTH�"� `�P�#�����S�
BETO)F�0#SɦDn�w�x�.�UNy���91���2}!L�8  � �0���B���@������BISPp0E�RIC@�A)$F�SB� ��CURR �Bm4�!�dbg.���������0
`U!R�E}pd0W0������ NEW��2�PPIP�1_P9Oa�EK_Ӏ_R>��E_DBG`���Tp���3��4��5_QޕsEOTF7 � $��P�$�`x*�nfpNCi ?�cJ�f?�*dJ�*g ?�7fJ�7i?�FdJ�Fg0��Td��TfUP��9 ލAEPCR7A�� ��ل� L�Hr  ��%�4��00��2�X��0À3KIPTHE�RJ�ـ���KEf��0�&��WV�2��Eð;0�0��PHK-1��@��� RM��CH�S�PTL�0�$H�z�SW��BBONLC�$B��2pfbgF"WF �1t��q�zE"�!� s_W;6�AND1o�\�!ND2v3v�aS� �A� ����M~�� | $�0 �@g�e�*f�7b��Ff�TfADAP�!�LG�CSENS�Y�r ��EVP�!�� 4?p�Oֱ o3�$F�r�r7cr Fa�Tarm�'��&�{�&�!4�&5�&6�"��f��ʿܼ�� ��B��6B�6��46 ��65đ͒0�7w�����Pe@�V���TAI����)�A3T��	TX1�'EP>���\GP�0S��$��\O OVӀI��"[�AM!ܒK5M� AF��^1BEF֦LNd]�+ù�%@��� mq `�ePPW)��:3�6i r��TRK�:�1�9MANU�qZ2m�D@D��AASR�EA � 	�y�&�`��  Ր�7y�q1^0Y6>H^1MIDU��If�!�����`�+�DEQ�w�CD0�!je�O �>P 4 ^'�q l&�S�������Q!�&P $ $E�LE�caQ�q5Ԇt	S���C����<;��r:�{:�0�TVPK �P� UU�uR�:�MU �eY�U��T� ���S$��S6XS��R���W������FW8�dBd��LAR�*�e *�)eO$`�O$p�O$��ЁQ_7�gUSh���cEC������PW{���_Og�#�e �f �eu)f��bw|�t���DI$񲄵@Ewr~pLEw@|SIZ5RxVu�D��BOAR�C@h� ��� `��a p��r{a�r�Q�U$VENDր���OEVIC1xD D�#j~�JւV}�IN�`�t�1��q;�MA0�CwpFIB�URf�f�~,E p $,B�/�,B/2��F,�O���,BC��Ǳ��TO�ԩ�_R.@M�����މ$BUP�� 4 Аo�-����p��?!L��!�PU�RA�PREFLO]W�OSTi�Rwp�+���A�0�������&��S_DlqdM�ఽ�T��d'���MF ST/@���n��t M�A�Ԡf��ر�$���΂qADJD��#NE�Xc���4���T_P�!h��1M�b�#( �Æ8�S_!���$�HaO�!�,�PFL� GAP�2I� �����BJWT`�C�Y�p�x���[�!�9 $B.s !r�@�-TOT�@�U�!rU�IApT�WAR~0DV���Ahz��r�Y^v��<�KG?r��0�k��"XsNp  �$ASCFl�"( ��O���#^��c�Qc�?!*�W�GLO�BЯ"���� NO-T�!$��IC9!�!AV��Y�\�$�"�5�1p��W_S+HF[W$1X#Ɛ"�I-�\� ?�t�RY��3`���p�3P�L@M��t���E�F UIF�o�0�O|p��!AD���\�APCOU9P����# @��(��-�
 5�x�EQ:{��@MMY��T����T���
P�0US�TOz��  ���{P}�� 
D;UE�EMG� �A7% ,QMG��� ��NOѠR�֨�7������& ! ����э����s �2T-�IR2T�q��)E�p�X`M��?��MI�T�CTSK_�WAIII��VG�	� S����7���T_GBUF����g�C`�ABNe��`������������D>�=����GcSIN���REd���1CT��NX�­�L�p�7���SA9VH��_PD��Iњe�W� LTn���PcIP�s�0BGa` ��[џ�fџ�qџ��P�"@��SPC�'� ,>#���b�A� ����� ���PPA`z�����i2P��>�cHE�@i�?!k! k�r��bk�"j�� �"`�B���Sp�B�R�B�����_FkIL�W�pBUN�0〷�b��F_��.�<�0wp��N�PSV�O �C�0a��PR>DIO�И�s��p��TMB�^
P�AP��� ��_'DYNe1i�Wr�F.�`KEYe0G��`@8�BF�1�@��� l$#�RPR�OU,$�C"� �B@bCAL��@`�`T��i�P��_#!RTy#H��0A��� �$$CL�ASS  �����! � �  � <0S�A�'�  ㆹ!I�RTU�0�/� AWCAO���A��3� ��!�!EAɐ s2�(0504;52�!?�Q338 b51:5J5J6�?�?�? �?�?�?�?OO,O;96EXE<
01?C? U?g?y?�O�O�O�O
_�_._@_R_d_?OɐS R!>gA�%�_�_ �_�_�_oo'o9oKo`]ooo�o�o�o��3�NLG 2"< ��q_qC?lK<�!A���okK�; �Bд!J X5� 2��%�c��General Purpose� �MIG (V�olts, t�)�p\ ��p
AW�MGENL.VR��vA*EGLM#G1�x�C1
�rB nu�Pxv�g�q�!�}<��N�`�r���sF�o�hC�NV 2	"<�2���sG 4���$���� W�6�{���l���ß�� ���؟�/��S�e� �����z���ѯ���� ��+�=��a�sL� =�����C�ܿ�Ϳ� $��H�Z�9�~ϐ�o� ���ϝ����ϣ� �2� �V�h�Gߌ�k�}��� ������w����@�R� ��v��g������ �������	�N�%�;� ��_�u����������� &J\;�� �gq����� F%V|[�� ����//�B/ T/3/x/�/i/�/�/�/ �/�/�/?,?��J? t?�/�?�?�?�?�?�? OO�?:OLO+OpO�O Y?�O�O_O�O�O�O_ $__H_'_9_~_]_�_��_bNVWP 2�&��\�dT 
�_oo0od}UST�OM 2&�l  ;o�o�o�o|�	�d�enrDEFmSVpR&���P�<�o�sDefault Sch A*wN`�� �����+��� a�s�J�y��������R�FBKLOG1 �@[mTlaBG������#�5�;�ۈ2<���C�  s���𗟩���ۄLG_C�NT  [moa��RIOEX 26[lDEeA Ec���	�@=i@=oa�a�
Weld S�pee�a�cIPM  �f�x����������ү���Eb �$?���none=k�#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q���������������R� 2��\
��@"��13-AUG-�23 17:36�:56�A23�0813Ee1�736�Eb̐��Q)	Undef�inO�����
F0���^����;��A>�?��W��m����� %
LAB�_L�D_1=j@Ed�ac^�@ig���Eb
�oB�����:��
������ ���������1! 3EW�{1/O/t/ o/�/��/�//>�/T�/?�@)?C??g?�/���? %�?�?�? �?�?OO+O=OOOaO sO�O�Oz?P?�O ?�O _�O'_�O�?�?o_�_ �_�_�_�_�_�_�_o #o5oGoYo<__�o�O �o�o�o�oloN_`_1 CUgy���� ���	���o�oB� �ou���V���.�" ���)�;�M�_�q����������˟ݟ+���B�OTF 2
T�?����:�Տ^�xp�G�a�=���*�@�󭯿�I�PC�R 2�p�!B�H��*B���.��C����!�ffA��  =�+{B�P5MܠT�"��Ԁ�W�OܠT�#����������	����2345678901���5�G�Y����à���@��$�@����C��޵<!��:#h�SR?AMP 2��:!�$���2<7Y�RGSEL R��   	�Process ,�1��2|/9�P*T��8�4a�t�5a����`+����*J��8a���ܠT�_� �*A|�v��A@*�B�&��<!�Ѭ�Vol�tag�	v�s�a�<�DwF�X�@]�ylس�h��Wire fee�d sp����IPMa�<��M�a���  ��a�����*�<� N�`�r����������� ������D��z�  �#��E� B�<!��o���ݵt��V���ѓ�Curren=t�Amp� ua���?Q-? Qcu����� ��//��h!��h% h!��h!��h!��h!�h!�,�/q������� ��!���!���!���!Ґ�L�/8��?�����Z�� )h/�	K/�?�?�?�?�?�
��S R&�$�A�4ᨵ!O3OEM�? �:EO�O�OSOeOwO�O �O�O�O�O;_M___ +_�_�_a_s_�_�_o �_�_�_Io[oo'o9o �o�o�o�o�o�o! �o�o'i{5G� ������/�� ��w���������я �����+��9M�k� a�k�}���)�ß���
�������,9բ�UPܠ ୔=��o?�33:�>>7�=L��>;�,�U!��"��#��$��Lf�X'�K���?^�r��>��r� ?J2�`�WIRE 2!��<������>��3�>�G(=��J*]�SCFG "��v��#��|��������O���#�OU�PLҠ#��� j�,�����w>��w;ۿ O���_��ѿR�I�[�>��NB  `%��� �USTOM �$�
6c�ɿ �E�MGOFF %l�6�#�LO*��&�ϑ'A��P�BM� �|uf�x  ���
,<�����a$��f�~��PCR ' �&~�@�bD�CE�5 �����D�_%��M�5 p���%��