��   	��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����AW_SCH�_T   � �$CMD_VOLTS  6�WF?AMP?P�KU
FREQYU�LSE@SPEE�D@TIM�FD�BK:�UOMM�ENT ���$$CLASS  ���������� VER�SION��  ��I�RTUAL��A�WE*  R �� t $ �<A�  +��?���F�����F Xj|����� ��//0/B/T/f/ x/�/�/�/�/�/�/�/ ??,?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�O �O�O�O�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o �o
.@Rdv �������� �*�<�N�`�r��������Runinx����م=��ͩ��	 Burnba�ck��
��  Wiresti2���@����ٍe� OnTheFly?�