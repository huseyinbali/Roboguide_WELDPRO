��   ��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	TO/GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1� � �CLo:o � �AX{ � $PS_�T�I���TIME� �J� _CMYD��"FB�VA >�&CL_OV�� oFRMZ�$DE�DX�$NA� =%�CURL�qW���TCK�%��FMSV>�M_LIF	���'83:c$�-9_09:_��=�%3d6W�� �"�PCCOM,��FB� M�0�oMAL_�ECI��P:!o"DTY�kR_|"�5:#�1E�ND�4��o1� l5M� %��PL� W ��  $STA:#T�RQ_M��� K$NiFS� uHYsJ� *hGI�JI�JI�E#�3AZCaB�A� ��$�ASS> �S���A�����@�VERSI� �G�  �~QIRTUAL�O�QS 1X� ���9@ ��x_c_�_�_�_�_�_ �_�_ojP5fBe&m� Q^oLm�%9�m��*��pg����7�t�� �ۄKo�ooql�o�o �o$�kW]r@F������d�������=L����8�?�9���@� Y�~�������Ə؏����� �2�D�� �1Uo�}�g����D  2�Ο�����(� :�L�^�p���<���� ����Я�����*�@<�N�`���2P��(� �������ܿǿ �� ��6�!�Z�E�~�iϢ�؍ϲ����$4 1�N\���L�k�cM��K�&�IOQ�RL�m��L���A�+@�xr@w��h<8	�<�?k(<$�4��k� \ߵ��ϕ߀߹�T�f� ���ߤ�1��U�@��y���Wzr�Wi-t���� ���p���l�����1�C���%��345?678901c�k� ��񍟨��������� ��`�"4��
�� d���v��� �J�*N<r �����\� //8/��q/�� �/"/�/�/�/�/T/%? 7?�/�/j?X?�?|?�? �??�?>?P?�?�?O TOBOxO�?�?�OOO �ObO_�O_>_�Oe_ w_�O,_�_�_�_�_�_ oZ_+o~_�_
o�_^o �o�o�oo o�oDoVo $�oH6X~�o� �
l����2� D��k���J���� ԏ��N�`�1����� d�⏈�v������� ��J���*��N�<�r� ��ڟ�������\�ޯ ��8�����q�į֯ ��"�ȿ��ؿ��T�%� 7ϊ��j�Xώ�|ϲ� �����>�P��Ϝ�� T�B�xߊۙ��ϱ�ݎ,��(����U���$PLCL_GR�P 1o��� p(�?�  "�4�,�W�(�{� f������������ ��A�(�2�t�