��   �A��*SYST�EM*��V9.1�0214 8/�21/2020 A   �����
�WVAMP�_T   �$X1  �$X2AY@�?�/FC5  �$2ENBA $DT  / �_R2 d E�NABLEDnSCHD_NUMA � xCFG5�� $GRO�UP�$z ACC�EL@�G$MAX_FREQ�z2 L�DWEL��DEBUG�PRwEWSOUT�>PULSEA�SHIFt 7TY�P4$USE_�AEF} 4$G{DO�  f0 r?�Np�WEAVE_TS�K �V�_G�P�SUPPOR�T_CFnCNV�T_DONE �p }k}GRP G2r�� _� ��$� TIME�1�o$2'EX�T� (1#&(MODoE_SW�CO3 OSWIT � U/ �PHAX6  4� � ECC$�TERMNnOPEAKno!AL  \ � Z�!I�$�!N_{VSTAR�#`!r"��"�%��CYCL42 Q
��/ � Tv"b �$CUR_RE�L_� �!3WPR�5 � 
$C�EN� _RI3R�ADIU�X�Iz ] ZIM�UTi!$ELE?VATIONg5� �N�CONTIN�UOe2q �MEXAC=PE�S��6  H~ �UE�NCYA�ITUyD4�2RIGHC��2LEBL_AN�G1 �OTF�_� 	� c $3A�bET���n3C!$wORGjHFBKjH���P��C��DLKDW�HR�E�_�3 �B�C��D�B�C�@�D�A�CCHG�G	Q�Fp	Q�F	Q�FINC�G =Q�F=Q�F=Q�F�AVC6PYC� _T�\#0�Y~P#�@SY��9H)@�UPD"0n��$$CLAS�S  �����Q��8 �P�PVER�S�1�W � ��QIRT�UAL�_�Q0 2��X� � {?��@�  Ha Dae�TWoio{o�o�o�`)dN 2 3k� Hf��uHe@O�Hi�oNc)a� � e� E`��i ��Ca��d �`z����=�����4s ����jpYq��w�r��1��x at��ujp`��i.�5t8q�q2�b�t���
�<q`����� Ca����̏ҏ�����)a�  23k
{TDaSI�L8� �����0h�?m�'����l�D� ����Ca��l����k�� � �2�D�V�h�z��l�FIGURE 8��o�v�Ha l�f��������M� (�H��󈯎�����Ŀ�ֿ�TCIR1��Pd�}�0�~�`h�z�D�Z�l���0� v˜�~����� ��$�n�jN� 2��4q�Ȓ���@��ʖD� M`g����������	��-�?�Q�c�u�`�� �q� �5)�ᐟN`���� ������˟���M�_��q������������k�Triangle��z�h߾�M ��Ɵ�ύ����`��/ L� &��g�n� ��	//-/?/Q/c/ u/�}DVhz��/ �/��9?K?]?o?�? �?�?�?�?��Lu�� Oe��O2ODOVOhO zO�O�O�O�O�O�O�O 
__.[�?._O"O�_ �_�_�_�_�_�_oo�&o8oJo\ono�mSC�HEXTENB � =��ctSTA�TE 2�k �|o�o�o �gWPR 7�6�L}�D�-�_OTF 		8��@)0�q�q�0��v)��uAȫs�u�@�  <#�
��?����mu_GP; 2w| ��� d�v����я㏡+