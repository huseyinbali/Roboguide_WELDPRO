��  	G��A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  .�pn�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@  �ALRM�_RECO" � � ALM�"EN5B���&ON�!� �MDG/ 0 �$DEBUG1PA�"d�$3AO� �."��!_IF�� � 
$ENA�BL@C#� P djC#U5K�!MA�hB �"�
� OG�|f 0CURR_D1:P $Q3LIN@S1�I4$C$AUSOd��APPINFO;EQ/ �L �A ?1�5/ �H �79EQUIP 2�0�NAM� ��2_�OVR�$VE�RSI� ��PC�OUPLE,  � $�!PPV1C�ES C G1�!o�ft A> �1	 �� $SOFT��T_IDBTO�TAL_EQ� �Q1]@NO`BU SP?I_INDE]uE�XBSCREENu_�4BSIG�0�O%KW@PK_�FI0	$T�HKY�GPANE�hD � DUMM�Y1d�D�!U4� Q!RG1R�
 � $TIT1d ��� 7Td7T� �7TP7T55V65V7*5V85V95W05W>W@�A7URWQ7UfW1pW1zW1�W1�W 6P~�!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$Nb_OPT�2� � �ELLSETUP�  `�0HO��0 PRZ1%{cM�ACRO�bREP	R�hD0D+t@��bl{�eHM MN�yB
1�0UTOB �U�0 �9DEVIC4ST	I�0�� P@13�r�`BQdf"VAL�#ISP_UNI��#p_DOv7IyFR_F�@K%D13�x;A�c�C_WA?t��a�zOFF_@N.�DEL�xLF0q8�A�qr?q�pF�C?�`�A�E�C#��s�ATB�t�
��WELDH2/�0 =s�q"QING�0$�QA7P<D2�4%$ASd3�B�El�P�_��BUC�C_AS�BFAI�L��DSB��FA�L0��ABN@��NRDY���`��z��;YN��SCH���pDE���yp�����8���|�STK>���	���	�NOj�?�ڂL��d�U* G���9  ���������߇Ɨ�Ɨ��ԘS_FәE���F�ƗSSŘ��P̂1 �ON�F�HO�U�D�MI�1�D�SEC`B�y�i �HEK0~��G#AP������I� � gGTH���0D_ȡ����T= ��륌�
� �p}�9!K���9!Ɨ�UN14��5��#MyO� �sE � �[M�s��t�RE�V�B��������AXI� g�R 7 � OD}`��'i�`M�m�� ����/�"��� Pŵ�eaX�@Dd� p E RD�_E���$FS�SB�&W`KB!�EF2uAG� J��  "��S�� V�t:5`��QC,2��a_ED|u � � C2��f�S�pa�l �t'$OP�@QB�q���_OK"�آTP_�C� ���da�U �`LACm�^��J�� FqOCOMM� K�D�ƀр@�p���OR�BIGALLOW�� (K\��@V�ARw�d!�A}!��BL[@S � ,�KJq��H`S�pZ@M�_O]�՗�C�Fd X�0GR�@��M�NFLI���;@Uɠ�84��"� SWI�&"AX_No`����9���G� �0WA�RNMxp�d4�%`Lp�Tb;�� COR-�rFLTRY�T�RAT T�`� o$ACC@�TB� |��r$ORI��.&�RT�`_SF\g��CHGV0I�E��T��PA�I���T�e`5��� � �#@a"���HDRՃ7�2�BJP; �CO�I�3J�4J�U5J�6J�7J�8J��9��Ȱx@�2 ]@� TRQ��$%fh������_U����� COc <� ����
�3�2��LLEC��o�MULTIV4�"fѱAv
2FS�ILD��
1;�Oz@T_1b � 4� STY 2�bv�=��)2_�p�:��� |9 $�.pڰx�I`�L* �TOF �sE�	EXT3ء�B3��22�0��@�	1b.'.�}!9�
���  �"�� /%�a�g�?s���!��;AآM��`Q  �T}RE� " L�0��	�`��pA�$JOB��E����$;IG� # d�,/ >/P(���#��ނ_MORc$ et�F͠�CNG�A�TBA �6c� :/�9��0�19@�G;P/pH5��?�%L����Bq�1��&rJ��_R������;QJ@��8�<J� D81 ��9Q��2�@��:�}Rd&� 
�	�rG�R�`HwANC?$LGw� �a2q�͠�Z�/���
0�2�R��Li�0�D��)�CDB`�C3RA�c�CAZ�`�H�ELT��FCT<�.�F"�`�)M#@�AI([O(X� ���
1�Rw�w 3�/�S���1��5�MP������HK&AEGS_SH�Q�W�ЅN0S��Z����'/  v@I#�Aq��Rc(��STD_�C�t�Q�3"US�T�U��)kTI�T�a~Ф	%�1IOy���@_Up�q���* \����UpOR@zs`b��}�~p�`O~@N�SYR�G`�q�e�Up�Љ�� ��U�PG`PXWORKz��+r $SK��l<�p1DB�TR�p_ , ��0A��0�c�B��W�DJDS �_Cd�`�sDPwP�Lzq�ё�s��DM�<wY����2��H�9N�p� Eb�A��-�bHaPRi�M�
�
�D�� ��. �q��1$�$-ZB�L�y/�������0���;�P� 1��t�ENE��� 2����a��v��r3�H $C��.$L`�/$�s���t�w�INEV�a_D}�m�RO3���I;��~!�`�:���RE�TURN��2MM�Rj"U琋�CʠN�EWMA`#�SIGeN��AJ@#�LA<�|!�&P0$Po �1$P�@�24�M�;�O��S����a�o��v�Q�V�GO_AWT #�`�@`�>�QW�DC)�o�KCY� 4'"�1�(�����Ĕ2��2̖N�a���C�4��DEV�I�� 5 P �$��RBU��P�I̗P��3�I_B�Y�;�J�T�1�H�NDG�q6 Hv�c&�E�g㸣�#@�㗣͖�`���L��7w��`�Ѭ�FBڬ(�FE�����͔(��@�ܱ8� �МQ��@�MCS4�Ƞ�d(H����RHPWF��5�:�J n���SLA�V.�9�INP���J��Ш����:P +B�S6@`�`� B�� 1�FI(b��	��5OaQ'Oa9W	�NTV䲹V��SKI�CT�E*�@��b�]�QJ�_S�R_���SAqFv�5���_SV2�EXCLUv`J-�D~`L���Y�<{�HI_VRP�RPPLY4px���u��۶��_ML�v`?$VRFY_s�M�IOC\�%C!_>PS�T�]�O/��ţLSр��nt4Fq$y�͓� �`P�en�l��K�AUNF�����͕���ZqCH�D�$������ AF�� CPU#��TFq8ĳ?Pס ;4��`qT��c�� ��9N�� <��8@�TЀ�� ��g�óSkGN=�0
$U0 ������Б� *0e �b��b��ANNUN�����͕U0�4v`'�w ����>P���V��EF�`I�>���$F��&d`0OT ��nt��prTq��kqZ)�M��NI�r?'"�|�G~�Aޱ��DA=YecLOAD�ct�u�os5v�EFF_WAXIɢ@4�Yq�SO���s�`_RT;RQ�A Dy�Q�� Qt` E���� @�P�WP|  ��AMPC@E�� B�XT0]2Xl�8FDU�8E]��bCAB�C8�f*�NSj9PID�!CWRBU�A:PV%��V_T  �@�DI�%0cD� 1$-V�SE�T�2]3��1�o�
Fp]2�1E�_��lVEP	0SWAQ�0� 3d  A_0��OHfqPPAmIRAa]2B�`�n��� ��S��@�@�%��� C�P ��R7QDW�MS�P%�AXt/lLIFAEp�. uq:"NA! M2J%��?#M2C����-C�P��N�$ǁ��&��OV��V&HE���]2SUP�!��D:"p_�$��y!_:3(�%���'Z�*W�*�Q`�'S�ሢ�RXZ�@��qY2=8C��T��`��	N?���J�%Q �_�@� x�`I@�TE `��CACHt��3SCIZp&� ��%�NZ�oUFFI� � p��ct��os6wry�M�P%DF 8��K�EYIMAG�TM���C#A��F��Ɓ>x�OCVIEK�a�G�R�@LCĐ� �?�� 	#�D?P�4H� b�STo�! �BFp�DTp�D��D��>�@EMAIL��x�����FAUL�r�I�R���cPCOU��PFA�`TO��QJO< $�C5�ST v� IT��BUF�7� ��7
�4`*`� B*T5�C�����BAcPSAVuU7R \2:�U�W����P|T5�R��L��_*P[U���YOT���`��P2�\p�Z�?��WAXec+�=�XX*P�éS_GA#
� �YN_���K <�� D0�!p���M��� T��FƀY$݀��DI �E�`HO�P��aL����GKQF�&�㌁�a������	�M�\��a�C�SC_��K���`���d��RA�e�H�aD�SP3F�bPC*{I�M�S!sGq��a� U`�g� ��"��@IPD�0�c{0 tTH[0��dr��T��!sHS�c�sBSCQ�j0*�V�ְ�z�p!c�tf���NV��G ��t[0v*P	FAB`ds}`aǁ�SC�&��cMER|��bqFBCMP��v�`ET�� NBFU� DUP���22��CDy�p�P�C�G�ЀNO�х�O� �������PN�Cj�υR�@b��A���P��PH *ρL۰����Q L����o�B��@�j�@���@���@��1@�7
=�8=�9=�A ?�I�U1V�1c�1p�1}�U1��1��1��1���2��2I�V�2c�2�p�2}�2��2��2���2��3��3I�3TV�c�3p�3}�3��U3��3��3��4��N�AEXT���QTb ��Y`m&Y`:�d`����"�FDR�RT
PV���R:"ɱ\�r:"REM#FU�NOVM�c�A��oTROV��DT�P6�MX'�IN��� ���IND6�
bȎ`B`W`G*a�!�ȁ@J%0D!�RI�V�n"GEAR��aIO'K�lN }`����%(L�?@� m�Z_MCM50:! ��F� UR{�S y,́MQ? � �\p?4�@?4�Et�<�H�gQX����T�0�Pa� R�I���07SETUP?2_ U ��6S#TD�px5TT��L�p�לչ�7RBACNbGV T��7R�d)�j�%<��x`�IFI��x`X�)�A ��PT�M�AFLUI~D�W �{ `H PUR �`Q�"�R�a�p-P��$ Iܴ$p�S$�k?x|�J�`CO�P��SVRTl�G�x$�SHO#���CAS�S�p�Qp%�p��BG_������c���p�<��}�FORCy�-�DATA��X�BF%U�1�b"�2�a���/�[0��Y |r�N;AV`�p�����S�Bn#$VgISI��vbSCd�SEZм�V��O
���B�I� ���$POt�I���FMR2��Z Ȳ��1bɱ �`��ͷ��������@��_����$I#T_ᛄ"M�ƲϾ��DGCLF�D7GDY�LDLѐ�!5R&��J$~�M���C�[G@;	 T�sFS�PD\ Pz���cB`$EX_.1`��"53P5P�G�q��g] �L�x�SW^U}O�DEBUG��L��GR��4@U?��BKUJ�O1� O PO ���j���M��LOO,c�SMK E�R�A�T�� _E ^ �7@�� �TER�M %_)&�0ORI�a% `)%��SM_�`��% a)%��h(�b)%���UP>UBc� -S���^p�7#� _��G��*� ELTO�A�b�FIG�2�a��,@N$�$`$UFR�b$À�!0̖�V OT7�TA��pɰ13NST�`P�AT�q�0G2PTH	Jn���E�@�R���"ART�P�%�@�Q�BΆaREL�:9aSHCFT�r�aM1{8_��QRw���f& q $�'��0bvʰ��\s9bSSHI�0sU9� �QAYLOvp2aHa1��]в�M1B�ׅ�pERVH�Af��8l�-7�`��2��sE��RC<\�ׅASYM{aׅF�aWJ�'l�h�El�w1�If◁U�D�`Ha{5� gF�5PZs5@
���6OR�`M��Tw!��d��L0�01a�HO���e� �S1��OC��!��$OaP���a.����$��`䰚PR�9a�OU�sM3eV�R�K5�U�X�1��e$P�WR��IM�UIBR�_�Sp4r�g `3�aUDlӳ3SV	�eQ�d]f��$H�e!f`�ADDR��H!G O2atamaj��`���g Hz�SE������e�ec��ep�SE�?��i�HS����gh $��P_Dq�x����bPRM_R�}�HTTP_�H�i (��OB�J��mb��$��L�E>3cP)q�j �s |�b�AB_c��T#{rSYP�s@�K�RLiHITCOU�t���P��P{r��`l��P�PSSg��;�JQUERY_�FLA�!b�B_W�EBSOC���HQW���!�k�`�@�INCPUdr�O :��qH�Q��dR��dR�~p� �IOLN�җl 8z�R��d��$SL��$INoPUT_!$�Pڡ�P�� |�SL]A� m�����مՄ�C���B�aIO^pF_AS�n�Ї$L��Ow���1 ��"b�!I������@�HY��X�1�n��U;OP�o `�v����F�H�F�O����PP &c�P����O�ǒ��h�ru�M�A6�p l6� CTA0BVpA��T�I���E&P ��0PmS�BU IDC  �r��?��P>���:�&?0qЂ��+��⩀N�� ���IR�CAڰ�� r ��myԀCY�`EA@�͡��ҬF�&c��k�Rg0�AA��ADA�Y_G�B�NTVA�E�V�.�Ȃk5:�.�S3CA*@.�CL��G�"���G���6�sr���Xl2����N_�PC���G��7�tЂ�S ޱ��JrG�>�p"�� 2se����6��u���Jr�LABp?13� 9�UNI�9'�Q ITY���$xe�R���vЂM��R_URLT��$AL��EN�n�s�tg �Tv�T_Uk�� �J9�6�w X �����E��9�R����"] A�Ӂ��Jv���#FL9k���
Ӻ�
�UJR��x �mpFA�7��7<ҽD{�$J7��O^�B$J8g�7PH!�p҂�78�c�8���f�APHI� Q�qӶ�D+J7J8�����L_KEd� � �Kt�LM��� y <��X�R�G�ţWATCH_VA��5@~�Fv_FIELDhey��L�ҁ�z R 51V>@¦K�CT��W�
�r�:�LG��{�� !��LG_SIZut���� �����FD��I������ ��" ���S����  ������" ��A8�� ��_CM#3`���g�-F�An�����r�T(���2�ိ�� ��������I��������" ����RyS�\0  (�SLN[р|���p �@ڂ��,��s:rYPLC9DAU_�EApt�|Tuk GqH}R�a �BOO�a?}� C7� `�IT�s�03�RE��SCR��s8��DI2�S0RGI"$D���+��TH�t �S[s�W�� �N+�JGMTMgNCH� �FN��bWK}��{UF���0�FWD�HL.�STP�V�Q X�� �RS�HP�(�C�4��B+�=P0T)Uq�/��>�a�@��Gm�0PO��'���i�sOC�EX'�TUI{I��ĳɠ��4	1�E3yd��0G���	�c���0�NO6AcNA ��QD�AI9�8ttt��EDCS��c��3�c�2O�8O�7S���2�8S�8IGN��G���zm��43DEOa5$LL�A{�HAT��~F�u�T��$��l�B�ä���-A\aF��P��PM�p}� 1�E2�E�3�Av��!�0 �m{Qk3������?�=Q�u� ����FST��Rv Ys�R0P� $E$VC $[[�p3VFV �`�$ L4�F��P[�`=�[����Q$eENp�$d%6�_ ���q�q`�� �S ��MC-� ��9�CLDP����TRQLI]���	i�TFLGR�P�a+cr�1D:�+g%�LD+ed+eORG��/!>bU�?RESERVU��d��c�d�b�T�c� �� 	e/%d+eS�V 	`�	na�d>�fRCLMC�d�o�oyw��a*d�M�p��Ѕ��$DEBUGMASI���	�Q�uTu05�E���TQ�MFR�Q��� � ~��HRS_RUہ��Q�A�T%FR3EQ��Q$%0��OVER-���o��F�A�P�EFIN�!%�Q�]q[��s�dǇ \���q��$9U�@޲?�`G�SPS�@��	�sC~ ��c�W�sU��bq�?( 	v�MIS�C.Ո d6�AR5Q��	��TBN�c ��&1ˈAX�R���·�EXCESH�ºQ��M���щm�a���T�R��SC�@� � H۱_�����S�����PJ;PT�ċ &�i�FI��MI��� � �Po�]^H RCT�Ns�ȖOҚAҚ��Ԑ�C��u�ԐUSED�w O�@TЏ�PX ����������^P)�/��+eR� �pSZ��B�_FR�`T��\�Z_��^�CO>� P
HqK�čA�h�cu�B_��LICTB�� QUIRE=#MEO��O��)�1�L�PM�Ŏ �P���hr⛣�b��NDK����Џ4+��9�D�x�GINA�DRCSM\�S��0ё��S#��%�PST�L�ѐ 4��LO�̐�DRI��EEX���ANGk2k��O[DA�u���5�=���MFm����v�I��RA�U&�( avSU�P�U��F �RIG}G� � ��` �S'���SG&�T�� Rn�P~�P��r��#mqPGW�TI/��@��r(�M\�Qr� t�+MD��I)�ƕ0��q�Hϰk��D�IA���ANSW�"�mA�!�D})�HqOR�b�`�Д ��U��VB��`k��_P��_Lp�ѕ ���@�C��Np+������P�� ����Pƴ�KEI"��-$qB�p��zPND2rz�a�2_TX�T�XTRA�31�%r�&��LOw ���$�G�&T�F�.�|�g��_�ڲRR2����� .W�[A�a d$CALIĀ�(�G�1��2�@RI�N���<$R��S�W0t��%sABC��D_Jഡk����_J3�
�1S�P��r�k�P�-�3P,���vPk�\�J%shl��b�aO.AIM%p�bCSKPj��> $qs��J~�bQ����p������İ_AZ�b�h���ELAg�qO�CMPҳ�aJ���R1T�q)Y�1�i�G�FȀ1�K40Y
ZW�SMG ���dJG��PSCL���SPH_�0Dp��`k�=��RTER���IS0��_�0�Q�aAS�b�DIn�23U��DF^P��LWVEL�	aIN�R0&_BAL�0k�.��l�Jx3LDMECHPB�%rP�IN� �q���@|҂�2�ҁsP_�� ����Hp�b?������DH�t3഑�v@$V��R��41$v �q�rV��$�a��Ro�����H �$B�EL �w�_ACCE4(�S'%qa ʐ)_� �q��TJ��C-*�EX�RL6��& c�w'��w'.�W)�'�m#�'36�RO
�_��A!"� 1�uu�W!_MG�sDD!1��rFW�`��]#=5m#X"�28DE[;PPABmN�'RO� EE2 �A�?	`��AOqO�X!�^P�_��bSP.�pCTR�4Y}03 Z�a yQYN��A���6����1Mwq�ѭr�0O ��CINC a�̱Z2A4˂:G��́ENC� L��k��!XX"Ʉ+�IN�BI6���E���NTEN�T23_�r�CL!O�r�@�pI�U� �Fj��\��@ia�yC��FMOSI&1�y���1�s�bPER�CH  k�q�  .Wұ9S���B�d��$��5)���A�"�UL �4��t����EF��J�V��FTRK��AY [�(�O��Q�"ecͰp/S�HB�pMOMcҀ˂O��`��T�Y3��0c�#�2��DU��7��S_BCKLSH_C�"�ewpV�p�3�j��caB�jA��CLALM�D}q>`��e�CHK�����GLRTY���ӁD��?�r��_�T_UMps�=vCps/1�Us�pLMT)�_L nt+�ywEs}�p�{rp�% �u�(>�aA�P�trXPC?QrXHI�۠%5�=uCMC7�/037C�N_��N6�4�t�S	FE!cYV�2��wG�p	��"x��CATD~SHþ�34iF?�xa�xFX�7�X�L "0PALDt8B_PCu'c_���� f"P��c&�uJ�A�T�a��?�'��TORQU�0/� Si�i0��R�i0��_W Ve�TU"!��#��#���I��I��I#F�尜�s�����+0VC"W 0�1Wd�1%�#089���+�JRK%�j�,]�u�DB� M��uНMP�_DL!�RGRV����#��#���H_^㈣� תCO1S�1 �LNl�� (�� 	�v 	�ۑE��3�����Z�V��M�Y����������T�HET0�ENK2a3#β#�CBӶkCB#C��AS�����۔�#�ӶSB8#$�޵GTS��1C0� �O�_Z�B�$DUp�W£�(5��DQnQ_�sjA+NE���!K$t;	��±AƵ����֥��LPH��§E��S(�@�3�@�B�� Q�j�T�q���V�V�� )�V8�VE�V�S�Va�Vo�V}�V��H�*�0�(ݭ�G�E�HS�Ha�Ho�H�}�H��O�O�OT��'�O8�OE�OS�UOa�Oo�O}�Oq��F���O�3�T��S�PBALANCE�_���LE;�H_ƵSP�$���3���>B�PFULC�������B��1�=U�TO_puT1T2	S"2N�a^"�@ 3�7a����"N#Ra�T�PO� `!��IN�SEG^"�AREV8X�@�ADIF�U��1���1��@O!B��a��dg2u��@�q��LCHWARL}2�2AB��feo��@��
AqXsX
aP�t)��� � 
p*��L!yEROB"P�CR�"l� ��CJ!_�T �� x $WEgIGH@i@$�d�)�IA�@IF�1N;0LAG�2�rS�2܃ �2BIL�OD�@`�@�STd �P��`�1 �������
]@J"�1� � 2��D�DEB�U�L� "~�M'MY9�%� N��m$�i@$D�!IQ$�W $���   ��DO_� A�� <�'& ���1��IB��N�C�(_�@��0"O�` �/� %\pT�@�A�[qT�O$� TICYK�� T1� %3��`(0N"P �#"PR��`�1�:5�F5� P�ROMPCE� $IRk��1p8�2�P�2MAI��2A4	B�5_��3� ta@R��COD,#sFU�0�ID_AP��5� {2��G_SU;FFې ��1�152DO=7x >5�=6GR��D[3 &D�1E�=Ev�D�$�6 ��H� _FIv+!9�CORD�3 �_"36�r�B|�1� $ZDT�5�m�  �%�4 =*�L_NA�!(0|�B:5DEF_I�H �B`6TF5�96$9602SF5@U`6IS��l� �!��94ySF3T�"]$4=��r"D �b��T,#Dh�O��"LOCKE��C:?L?0^7{QB@UME�B D2SD@UD�R&Bc %ES&DPT&B&{f{Q 1C� �1E�B1E2S1C�g�eH� P� iT� �uQ��� W�X�e�S�-��TE�a�$�� �LOMB�_r/w0�VIS���ITY�A$�O>�A_FRIWsF� SIuQYq��R%0H�w00�w3E#�W\x!Wh{��^vn�_�y;AEAS�;B5�Vtŀ��P�2�v4~y5~y6��ORMULA_�I���G�G� �h S.7e%COEFF_O1o r�$1C�G���S�~"�CA���/�#!GR��� � � �$�PF�"X� TM��W܄�U2�S���#E�R� T�T�D6 � M ��LL<D�PS�g_SV�TH�$v�6 �� G�6 � �΂SETUuSMEA�0�0��!�B��� � q�] g @����µ��Q��"�B(0�Q�Q�T��A�qFB�f1�P�Q��P����� �0RE�C�A���ASK_���� P�1_USER/�N�p? s�N�/VEL� N�? v�j��I�@� w�MT�!CFGD���  *0� ONORE�� ����� ��� 4 ����XYZ��C�@ J#�ʠ_ERR�� ����!��0���2!:����� BUFINDX��Ȣ�pR� H�CU��!_��1��A����A$Lt�OQ咻�@ ���GĂ� � $�SI;��p�0{R�V�O�����POBJE<����ADJU�"´FѰAY�AɳD���OU�@�_��1�B=^�Ta .�v�-��"DIR2�:�� ��ziDYN�ry�v�	T ��R^q� ��¿�OPWOR�� ��,� SYSsBU���SOP��H4�_���U�ˡ P�P����PAQ�����V�OP/@U�����)"f!�IMAGb$��&�"IMw��@�IN�p�?�RGOVRDk���R��P�>�i� �`�S�ՊL�PB�� ��P�MC_E�@4�[!N"��M��f!_"1d"�@�k�SL��E�� �^�OVSL�S�bGDEX�QNP �2g ��_k��a@l��@a@"�7�2�_"W�CZ��@�f�4�l�_ZE�R���҃�D�� �@נ��3O�@RI±D
��0�����ǡ�ܰLD��Z�T< ATUS��u!GC_TV�C��B�� ��Ṕ�Se!���@E�� D�!���s��v3�A?�$���XE@���\�p�;��㲠����UPPoQP!X�0.��]$3��7��PG�����$SUB��3]a�����JMPWAIT8��'�LOW�1���CVF�1+0bRK���&CCi��Rm�2_IGNR�_PL��DBTB2 PsQBW�0U2��U� TIG�j0=ITNLNS��R���R]pNj0��P�EED��	�HADCOW ��ʰE�p���PSPDD�� L�A'�P"�0UN���.��Rw�q�LY�@�  ���P��D���a$���f0� LE��� PA�P����yP�~�S�ARSIZ�4�@�CMQܰqO>@�9�ATT��p�-����MEM�"f!�TUX��}�qsPL�0��� $��~�aSWITCH	Z�!WͰAS���1"LLB~��_ $BA+�D�S�BAM��[Å)��w J5����"6|�&Y!_KNOW�4�"k�U�ADz(���-DQ��)PAYL#OA���`3_D�7T��7Z3L]aA���>PLCL_� !}�D2�!��Q4��_6Fi9C�?:��B4[�I?8R�?70��[4B�p�Jq��1_�JI1i���AND�/�
��4I2]1���qP�Lh AL_ �@= -���!��<pC�uD3E��J3�0�F� TU�PDC�K��rR�CO��_�ALPH CfCBE0��(� O2L ����>�� � �� ?WD_1:224D��ARc��H�E�F�C���TIA4Y5Y6�MOMq�S:S'Sh:S4S��B% ADSp^V'S^V4SPUB��R?T�U'S�U4R���@�G@��  r�M,2� ,&�A��� e$PIm���CZ�7i`�T'9iIkIkI+c@�T�\f��\f�����\Bg�Wª��HIG L#�&�f&\  K��f�c�h\�i\&SAMPk�d�t�gps&� �3 o� Fq��z�Ut��_v �@ny�@z�����P]u�q�b]uIN�|�p�c �x�{�t&�z�x�t�{^�GAMM�uS
�>��$GETW�@����D�D��
��IBt���I�$HI�!_[�D�z���E����1A������LW��̆ Ì�������B�f� AC�CHKyг�ڐUNI_�`����B �H�q�uY�RS��|VX��GC �$BH �1���I��RCH_DX�����G��LEv�Z���嘩H��}�� MSWFLVn�QSCR��10���SN�Wr3��:�|w��PnyN�]�PI�3A�VMETHO�}モ���AX���h�X� ���ERI���t3C�RB�5	D�a�@F4�q\s��ks��LĐq�OOP\q��0�kq��'APP��F�И04�U�@��sRTբ�O�0���a����T`1���T`஺+`���)�MG�ѳPc$SV~�PD�G� ����GRO� ��S_�SA�!��ū�NO�@C���D�b��O ?%?1h�o�W`�"_e,���CDOA_��  UvP��u�h��g��h0����H3 �A0 }M�U� � ^��YLc�1�w��S �2Q��b�(����1(��nӽ1_đC�Z�'M_WA��� �w����Mj ��d0��A�3)�	(����PM���R� � $�Y�m��W"�n�԰L !51"��D �D �D �4D{ ��N� d�C#����pXjO�C�qZp���P0 �T� ���M��W�T�f�xϊπ��P��ّ��A_��� |SA���:Y l�'Sl�4S�Z����-ZR!\�H� ��P�鲥�* 60P�P��PMON_QUp� � 8�QCsOU���`QTH� sHO[� HYS�3ES�" UE º�O5$�  ? P� �|�3�RUN_T�O���PO�b�P� P� `C��/����INDE��ROG�RA��' o�2��N�E_NO�`ITx�Q� D INFO��� ?!�
�m��v��OI�� (p�SLEQ�f��e� ʗCD S2���{ 4�ENABN�>^ PTION���ERVEdb[rac �3GCF<� @b J�Уqh�h��R�\n��PEwDIT��� �/�R��K�Q�c��E��sNU��AUT.��COPY�Q�`,ra:�M��N +*��PRUT�R "N�OUC�a$G�ep$��RGADJn��� hS@X_��AI͓���&���&W�(�P�(�&�c� �N^�0_CYCN�p/RGNS8�P��`�LGO7��`NYQ__FREQ�RW�p��f-1SIZK8�L�A��$1�!5S�p�eCcREo���8�IFa��NA q%k4_}G��STATUS�<��VMAILrbAx�1�LAST�1�aA�$ELEM<�� �9�FFEASII�KrD�t��2�� �F٢�pn�I� l��$2�a���KBAB$2�@E� �`V�1cF�BAS�BdEn��QU8�`�`'�${A�GRM�PREC�qؐ�C`���`��1�D � �2�S�[�	"B 2� �s���t V�BW�B�Њp�ѡB83W�WߔDOU�Ӕ�O��$Pݡ�@�G�RID�2BAR�S�gTYJ�2OT�O����� Q_"�4!� �RnTO��9�� � ����P�OR��S���SSReV�0)�T�VDI0�T_e``#dr`-g`�-g4+i5+i6+i7�+i8a�F?�<�~O $VALU~C��D@pF8��� !E;��S�1�۠ANõb�1�y�12ATOTAL�_�4I@rPW3I|vQ(tREGEN&z;r��X�Hu����f���TR�C�2&q_S��w;pأV�!��rsdBE�3ݠB`���cV_H�PDA8��p�pS_Y6����>6S�AR��2�� h"IG_SE��p�R�5_d �tC_�V$CMJ�C�T�KDEE��b�I:��ZS�-�N1�bENH�ANC� p��AG�2A3�qIN�T`�!��FZ��M�ASKʣ�@OVR ����ݠ��1��WV	 �byU�A�_'Fd{>�V�PSLG%��a� \ �?57���p�0S���4f�Us�V|��s��7a�UP�TE���@�' (cq��J3�.N3IL_MM4�VQB۠��TQ�𖣷R�@C����V�C-��P_�'�7�MN�V�1M�V1[�2j�2�[�3j�3[�4j�4 [�����ޣ�ޣ����;IN��VIB�'������2�2#�3*�3#�4�4#��� 6�O�2���D`�Q`�����PL�0TOR ��INƵ��R���L��T $�MC_F  5�B��L ����pM?�1I���OS ]���f���KEEP_H/NADD �!B�h@L�C�ᐐbĮQ�t�c�O��A� ���p�cë�c�REMz�@bĺ1�R�Ŷ���U�4�eb�HPWD  ;B�SBMӁ�P?COLLAB���`he�qq2� IT0��&"NO�FCAqLE����� ,���FLK��A$SY�N��`�M��C@��~�pUP_DLY��=�ODELA�л1ښ2Y��AD������QSKIPN$�� ��Pb Op���(���P_b ��� � ��� �׵ �s � D`��Q`��^`��k`���x`�څ`��9�!�JS2R� ���AX�@T'3���A�� >�p��>���RDC�a.T�� ��R�˸�R`1ɺȲ
TRG�E�4CгXRFLG����ŐSWX
TSsPC��!UM_��ؓ2TH2NRQ�k�� 1� �	���Q8 �� D� ��:�l@2_PC�#��S���A.0_L10_CL2����́ �� b�'` ����F(������� ��+U��г+� �b9�lCHЅ�����}�~DESIG��.'UVL1��1��Hvs10��_DS�h(�@��F  11�� l3�i���o�F&�AT��q$]Q07�'+$�  ������HOME�й2�������! �3�� DVhz��� �4������	/�/ ��5��>/P/b/t/�/�/36��/�/�/�/??S U�!7��8?@J?\?n?�?�?-'8��?�?�?�?�?O-%�S���  @�A�Pp6���E�T� T���D	v�C�IOՑ�IIp@5�OB�_OP�ESr�C޸POWE���# �@_п��"t� �Z�BR$DSBf�GNAOs�ЩCq�`�M����Z�CIk T_SP5E%�z�MD�W���Â�a��DBG_\@PU�����SEq<�̀ 2�4C=�ޤ2S232�E� Ɍ��7Eo���IC�EUSs�U�ARsIT�qqOPB.�ޭbFLOW�TR`�@r���P�aCUV` �aUXTҁ�a���ERFAC;d��Uv�`-"SCH��� t3����QH�@�3$�p�pOM����A�  t��UPD�����qPT�@Y�E�X��x�c!�FA��e�G��rfq � �цp�� (�AEL� �3u���:R�;�  2� ��S���@�	� ��$X��_�GRO�UQ�sT\ ��vD�SP�vJOGLIB�cF����,a7�N��Ф���ސ�fK�`_McIR�q�T�MT��AP��c�*�Z�`�SYq�t�]��@��BRKH�avl�A;XI~A  f�@��q��rρТu�BS�OC�v��N��DU�MMY16,�$�SV��DEQnSFSPD_OVR.�����D؂�sOR$�P@N���Fv����pOV�uSF�RUN���F8��a�soUFRAN�TOld�LCH�Ҥ��OVׄ8��pW- ��sy��P�����_8�� }@E�TINVE$P.KAOFSǐCSp��WD ��������R#��ÀTRO�R(�FyD��(�MB_C4��B� BL~���q0�6��qPV�adB�`� ���G1�D�AM�B�$��`r�����_M`H��b<��C��T$�����q~CT$HBKX�a/�ءIO_E�Q��PPA۪��������R��DVC_�PdCI�q`RI��D�a`�1h���`�3h�@��"��`�pׁUdC�p�FCAB��^B[�"��&�k�h�O�U�X/�SUBCPU_R�pS�����Z��`���I�Z�?R��$HW_C� t`����N��N@pNp�$�U-�z�t�m�AT�TRIEЁ��pCY�C��ұCA���F�LTR_2_FI�qCsY��fV��P�{CwHK_�`SCT�F_m�F_w� ҉��FSeQR�r�CHA�����A�Q�{b@�RS�D��bQ��s`QP_�To�? ���q`EM�@��Mn�T.��Np�.��Ӷ�DIAG~uRAILACV���MpLO��f񳆞<�$PS�r`B X�����PRJ�SZ�J& �C<�C 	���FUN��aRIN�Z�Y@��?�����S_�pu àh�@�Ѥh�-�ѤCBLCUR}��A�������DAx�i�����LD�`ˀ����qr� ���TI��}��Np$CE_RIYA��oRAF�P�SXG�[ L�T2��Cs̅�C�OI��DF�_L�@P��as`LM��SF;HRDYO,�ѐRG �Hb���Y@����MULSE�����Ǽ�s�$J��J����FAN�_ALMMWR=N!HARD`@�f�fs�2Vaz�R�_,��/�AUR�R3ԇb?TO_SBRU���p�
m�>�G�MPINF�������n�REG`FNV�`ԖSb�DPN�FL_Ž�$M�����cH��Np(/C�P�� ��b��PӐa�v�@$qA$Y�R��a	}r�S�7� �7�EG�@�s�ˀ�A�P�D��25p�����D�AXE�wwROB�zRED�v�WR�Pk�_���S�Yh��Ϡ&S!'WcRI�P�M�STOPP�s�`l��Eo��@"�6��f�pBa ��rh&7�ӝ�OTO�9�@Y�ARY�s�"0�ѝ��B�pFIM��s�$LINK��GkTH�"
pT_^#ʽ��8���!XY�Z�b�*9�&OFF�Ő�"�P� �(� B�p4�D4��mP�`E3FI��^7K�nSÄ4��t_J,aNr���#0��[ w$�*30��9`�Е1���2C#Q4�D�U�³�3%���TU�R X"�E�!�X0 `�7FL� l�̳P�$@5d)35�Ғ� 1��@K�pM /��6�������cORQ�ֺqn�8��
J�O N��E���q���DOVE�A�RM �`�Aj
Up
Uv	V�aWαWpTAN E��!
QL�Q�A�IP ��QU�AW�Up�UL.S�qER�qr�	 �!E��Dp��TAQNpa5`�ҫ'��׶��AX��Nr�ᝰV��" +e��7i��7i��6j� 6jq 6j� 6j� 6j06j1�06f��3i��Ci ��Si��ci��si���i ��i��i��i�a�ioDEBUE�$@�`L��tqڒ�"AB���ء ��CV͠D� 
�rq�r�u5��w�� �w���w��wq!�w�! �w�!�w1R��0L��".E3LAB[2�EA��N�GRO���2E��B_�ѸVM$��U0�� l����E��y��ANDr@ ��T���%�Qy� ��M^ �������� NT, ��+�VEL��eT5���=�줚E3NAc��� �$��ASS  �������� x�ʐS�I������㆔�I���������AAVM, K 2� �� �0  �5Ȋ�����%� %�	H�9�\����!�J���n���8������G������АB�SQ� 1���? <�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A�pS�e��L�MAX���Vh��5�  d�z�IN����y�PR_E_EXE����ȵ��D�����АIOgCNV*B�� ȑ��P���0��1��IO�_�� 1ݛP $͠�r�]��Z��?�h���}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c��z�LARMRECOV ������6LMDG �FQ k�LM_IF F��h�� "�4�F�T���wωϛ���Ͼ�, 
  ����b�n��1�C�T�$��x�_ߜ�[�����������s�NGT�OL  �� 	? A   >�P��z�PPINFO Ż Ķ���8����  �»� �者�����6� �2��l�V���z�������� ���(:L^�p�����غP�PLICATIO�N ?-�����Ar�cTool  �
V9.10P�/30O��
8�8340-F0S@105-">47DF1(��None��FRA� 6�p�_ACTIV�Ep�  �7�  ��UTOMOD� ��5��CHG�APONL$/ �8#OUPLED ;1�� u y/��/�/�CUREQw 1	�  T�)�,�,	�/	5� �4���"_ARC Wel���AW���"A�WTOPKS6HKY?���/�/�/?v? �?�?�?�?�?�? OO O*O<ONO`OrO�O�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xojo|o�o�o�o�o�o �o�o0BTf x������� ��,�>�P�b�t��� ������Ώ���� (�:�L�^�p���ܟ�� ��ʟ�� ��$�6� H�Z�l�~�د����Ư ����� �2�D�V� h�z�Կ����¿�� ��
��.�@�R�d�v� �ϚϬϾ������̹%�TO(�/#DO_CLEANE/�|��NM  -� �/������ ��.DSPDRYR��&V%HI" ��@��~� �������������� �2�D�V��MAX@� c��1T't�Xc��sp"s�PLUG�Gc d�p#%PRC*5�B����m�_����O��>��SEGF< ^0.7�߶߀~������1LAP[�n03 2 DVhz��������TOTAL|����USENU[ �h+ I�M/2� R�GDISPMMC�^021C+3�@I@�"h$OY�{�I��RG_STRIN�G 1
4+
��M- S�
~�!_ITEM1�&  n��/??%? 7?I?[?m??�?�?�? �?�?�?�?O!O3OEO�I/O SI�GNAL�%T�ryout mo{de�%Inp�@�Simulate�d�!Out�L�OVERRX� �= 100�"I?n cycl�E�!�Prog Ab�or�C�!�Dst�atus�D�@ce�ss Fault�\AlerT	HeartbeaS�gCHand BrokeZEWOY_k_}_��_�_�_�_�_�_ _��+_��/�_9oKo]o oo�o�o�o�o�o�o�o �o#5GYk}�_WOR: �+�q)o �����%�7�I� [�m��������Ǐُ�����!�3�PO �+1QY��{B�|����� ��ğ֟�����0� B�T�f�x���������үT�DEV\���p� �$�6�H�Z�l�~��� ����ƿؿ���� ��2�D�V�h�z�PALTm���{����� �����#�5�G�Y�k� }ߏߡ߳�����������GRIy��+E� ���m������� �������!�3�E�W��i�{�������3�+ R m��]���#5G Yk}����� ��1CU��PREG�Ύg �����/!/3/ E/W/i/{/�/�/�/�/��/�/�/[M�$AR�G_�pD ?	����<1��  	$�[F	[P8]P7��[Gq9/0SBN_CONFIGj@<;�A��B�1�1CII�_SAVE  �[D�1�3/0TCEL�LSETUP �<:%  OME�_IO[M[L%M�OV_H�0	OOR�EP��ZO%:UTO/BACK�1<9�2FRA:\{� eO{�0'`r�@{�H� �K��0 23�/08/13 15:18:50{r8{_-_Z_Q_�L��z_�_�_�_�_�_�_{��_)o;oMo_o qo�oo�o�o�o�o�o �o7I[m �������\!����  �A_}C�_\ATBCKCTL.TMH�`�r�p������oKINI����E�5�1z@MESSAG�0ρ�1D0ڋODE_D�0�6�5��O���wCPA�USm� !�<; ,,		�r0 <5q��e��������� ��������S�=�0w�a�s�����D�N�?TSK  T��O<��z@UPDT�͇�d��XWZD�_ENB̈́�:'�SCTA̅<1�.1WJ@�ODP�2<;�4W�)13-AUG-2P7:33P42O��@˿ݿ�1��F�L�ῠ߿*�7�`���
u�B���� ̐ � :�fϚ���j�R�OBGRPҨ�A�"�WEWE�Lp������6:5�6��D
LAB_"��_�D������9 k�f��nߟ߭���q�p����+4XIS�0�UN��Ԧ�1��� �	 I����Ck`� �	1! ��pګ{V��D�1�2���t��{V�Q��� �AN ���n� �$�)�Z��������0�3�MET��2�D鄰 PU�@n���@ �G@��6?�@f@,��@vo��>���>���='��?3^�>l��m?�&9�S�CRDCFG 1�<5�A ��� ��� );M�O{Q�9�� ������^ �?Qcu�� :'7}AGR=��2���C�NA#@;;	�}D�_EDˀ1�������%-I�EDT-���m/����@!~BI/:�r2p_FB/�/  ���%2�/6K�/F? 7��+??�/�/n?�/�#3�?'?OK?]>�?@KO�?�?:O�?�#4�O �?�OO]>�O_^OpO_�O�#5O_�O�_�O ]>x_�_*_<_�_`_�#6o�_ho�_]>Do�o �_o�o,o�#7�oWo 4{o]>{�o�oj��o�#8�[/ ��^=�G���6��B�#9��̏�^=����Z�l�����!CR�/"����X}r�ݟ�$�6�̟Z��% NO�_DEL��GE?_UNUSE���IGALLOW �1��   (�*SYSTE�M*L�	$SE�RV_��Lٗ�POoSREG��$£Lܗ�NUMŪ�ح�PMUC�L��LAYO�L��PMPALS��COYC10$�7�!�<%�]�ULSU�٭�9� ��Ls���B�OXORIɥCU�R_��حPMC�NV���10�M���T4DLIB�����	*PROG�RA��PG_cMI%�O�a�AL/Ŕn�X�a�B�ϗ��$FLUI_RE�SU=���ϯ����MR��������Wr?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q�������������%�7�I�[�6�L�AL_OUT ����#�WD_A�BOR>�g���IT�R_RTN  �Ā���NONS�TO �� O�CE_RIA_Id����0 � F?CFG *0���9_PA��GPw 1CUA�����C;���� ��C� C �� (� M�C8� @�� H�  CX� `�� h� p� x���� �� �� �� �`Rdv���?�{HE�ONFI�����G_P߰1C 1������/ /2/D/V/h/�KoPAUS��1��0 M�j/�/���/ �/�/�/?�/6?H?.? l?R?|?�?�?�?�?�?��?r,M��NFO �1��S  � 	�OO;�=@�B�B�QW��ڲ�B����jY�����B��CB���Õ���v2����IBB��L�A�D�B��jA{"�@^�@EC
�8O=�C�Ǹ�COL_LECT_=+F1��R�GEN/�����R�ANDE�C��GR��12�34567890�[W:ұ�SY_kV��
 %}�;�)�_�_�� �_�_o���_�_Too 1oCo�ogoyo�o�o�o �o�o,�o	t? Qc���������L��5V��2��K ]9RIOG !DYQ����`Ώ������TRr S2"�� ��
-���#��<��Y�_MORz�$w ��ŕ<Ařݟ˟�@�%����m{�%��%,�?���x�;СK��;ѷ� R=&��O������C4  �A����;�=A>{�Cz  B�${B�"  @Ңs��;�:dڍ�V�ARI=S'��?��z�(���/�d��To_DEFz� X��%J�������NUS�<��0��KEY_�TBL  �0�6B�	
��� !"#$%&'�()*+,-./�dW:;<=>?@�ABCe�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������h���͓���������������������������������耇���������������������9�p�b�LCK��	�b���STA����_AUTO_DO9��&�INDT���_T10�"�T2�o�V� TRL^d�LETE�����_SCREEN ��kcs�cU MMEN�U 1)�� < o�|�D�UE#�M��i� k������������ 6���l�C�U���y� ���������� ��	 V-?e�u�� ��
��R) ;�_q���� /��<//%/r/I/ [/�/�/�/�/�/�/�/ &?�/?5?n?E?W?�? {?�?�?�?�?�?"O�? OXO/OAO�OeOwO�O �O�O�O_�O�OB__��_MANUAL���DBc�j������DBG_ERRL�j�*�D� �Q_�_�_n�QNU/MLIM��[����
�QPXWORK 1+��__oqo��o�o�oS�DBTB_�� ,�]ģ�����o�DB_A�WAY�SD�GC;P ��=��1b�b�_AL`��b�RYЪ��ը��X_�P 1-��h�
No����|��f_ML�IS��
{@{��sONT�IM��������vGy
��\sMOT�NEND��[tRECORD 13�� ����G�O���u���
r��ŏ׏ 鏀�����<���`� r����1���)�ޟM� ��&�8�ӟ\�˟�� ���ȯگI���m� "���F�X�j�|�믠� �Ŀ3�����ύ� Bϱ�M�տ�ϜϮ��� /���S���w�,�>�P� b��φ�q�߼�+��� ���s�(���^��� ����=����K� � o�$�6�H�����~��� �������������  ��D��hz����bTOLEREN�CtB�QrpL��͈PCSS_CNSTCY 24?i%��P�Or�	 );Q_q��� ����//)/7/�I/[/�DEVIC�E 25�  �f�/�/�/�/�/??�,?>?P?b?��HN?DGD 6��`�Czu:O��LS 27�-t?�?�?O�O,O>OPOv?�PA?RAM 8hy8r�wUbD�5�5SLAV�E 9�=�7_C�FG :�ObCd�MC:\� L�%04d.CSV�aO"�c	_!�>A &6SCH>P�1�bN(I_~_�G�bFnR�Q�_�Y�Q�@JP���S�^"��a�>_C�RC_OUT �;�-�afO_NOC�OD�@<hw�MS�GN =^�G�#�M�16-�AUG-23 1�2:399P�Av`3�zf5:1�a�& Wzz�i�abN��`ra�M�����j��a�n�C�VERSION �ejV4.�2.11�{EFLOGIC 1>�/ 	�X�@Iy��QY}+rPROG_�ENB<��6ysUL�S�w �6+r_A�CCLIM�v���C��sWRSTJNT�F��A+q�MO�|�QPb�tINIT ?�
^��A� �vOPT�@ �?	6��
 	�R575bCc�7�4h�6i�7i�50��t��2i��X��%w>F�TO  R��ot�&vV�DEX�w�d�riP$�PAT�H AejA\��q����HCP_�CLNTID ?<	v�C �[Z�ß�IAG_GR�P 2D�I �> 	 @�K�@G�?����?l��>� �ٚ��8��ٜ5��� a�O�?��b�?> ��i�^�?�Vm?Sݘ�ٙf403 �67890123�45����� ��s��@nȴ�@i�#@d�/�@_�w@Z~��@U/@O��@I��@D(�XٚѠiQ@�6Tp6P,�� A�� � 9PB4ٜ� ٔR�iQ�
Т1��-@�)hs@$��@� bN@��@�ڠ��@�D@+2�	���-�2�A�2�P�R���@N@I��@D�@>�y�@9��@4��.�v�@(��@"�\��������пV��L�@Gl�@�BJ@<z�@}6ڠ0�`@*��$���@���&�8�J�\�V��=q@��F�@|�@33�@�R@-�?���?��`?�+�ϲ���������̑҂��-@_&�@�����!?�?� �,�>�P�b�t� V� �(�:��^�p��� D��������x�� ��6�H�&�l�~���� :���q�����ѡ��x������Y�̟�?�z���(�5�AF4� �?�L4R� (��@�p�8�Q�b@-: I �m@����%�Ah.�=H�9�=Ƨ�=�^5�=�v ��>{�(�=�,���,�^ �iQC�)�<(�U�R �4�����ٙA@hR?0���"��0 Vh4��t�8�����
/��>���y,"�R=����=��z<!(��7�G�T/G�(�8U 8U����(�$@9P��|*��uB�J����B�B��B%�(��T�/�.'�p5.�*11n,�\��=�-��cT+�a Bk B��BC�A��@�Z?؟�?iQ<�P�?�?�?�V �?O�?6O�+TOZB�ٙC�;
����$��9��4�B�ܻ��$O�O O�O�O�O��O�O#_2�>����>ˠ������>���@V�?j�_��'_u_��CT_CONFI�G EDo�c�eg�U�STB_F_TTS�w
�y��S p�s��V5`M�AU�p��rMSW_CF�PF��@��l�OCVIEW�PG'm3����?yo�o �o�o�o�oPrgo�o  2DV�oz�� ���c�
��.� @�R�d���������� Џ�q���*�<�N� `��������̟ޟ ���&�8�J�\�n� ��������ȯگ�|\KRC cH`��R!�� ��$�Y�H�}�l������ſdSBL_FA?ULT I�<h>߱GPMSK�W���PTDIAG iJ�Y�!�S��Q�UD1: 6�78901234A5O¬RC��W��Pb_ �ϝϯ���������	� �-�?�Q�c�u߇ߙ� ��j�?���
z���>�VTRECP(�:�
H�:�a���y�v�� ������������ *�<�N�`�r��������������=gUMP_?OPTION�P�F��TR b�S��PME�UY_T�EMP  ÈW�3BQ0m �L1WUNI`�Um��YN_BRK �KRo=fEDITO�R��F�_�E�NT 1L� � ,&	LAB?WELD_2��mL�&
� _? �(1AF���ֲ�������/ �;/"/_/q/X/�/|/ �/�/�/�/�/?�/? I?0?m?T?|?�?�?�? �?�?�?�?!OOEOWO��PEMGDI_STA�+am�R� �NCsC1M'k �����O�O��
��d ��_'_9_K_]_o_�_ �_�_�_�_�_�_�_o #o5oGoYoko}o�o& �o�o�o�o�iQ�o "4FXj|�� �������0� B�T�f�x��j�o���� ͏ߏ�o��'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uϏ�}ϫ� ���������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m�ϙϣ����}��� ���!�3�E�W�i�{� �������������� /ASe�� ������+ =Oas���� ���//'/9/K/ ]/o/��/�/�/�/� �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgO�/�O �O�O�O�/�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oyOko�o�o�o�O �O�o%7I[ m������ ��!�3�E�W�qo�o ������Ï�o���� �/�A�S�e�w����� ����џ�����+� =�O�ɏ{��������� Տ߯���'�9�K� ]�o���������ɿۿ ����#�5�G�Y�s� }Ϗϡϳ�ͯ������ ��1�C�U�g�yߋ� �߯���������	�� -�?�Q�k�Y���� �ϻ�������)�;� M�_�q����������� ����%7Ic� u���Y���� �!3EWi{ �������/ ///A/[mw/�/�/ �/��/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO e/oO�O�O�O�/�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCo]Ogoyo�o �o�O�o�o�o�o	 -?Qcu��� ������)�;� UoG�q������o�oˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�M�_�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� ��W�a�sυϗϱ��� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�O�Y�k� }��ϳ��������� ��1�C�U�g�y��� ������������	 -G�5cu��� ����); M_q����� ��//%/?Q[/ m//5/��/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O7/I/SOeOwO�O�/ �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'oAOKo ]ooo�o�O�o�o�o�o �o�o#5GYk }������� ��9oC�U�g�y��o ������ӏ���	�� -�?�Q�c�u������� ��ϟ����1�#� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���)�;�E�W�i�{� ���ϱ���������� �/�A�S�e�w߉ߛ� �߿���������3� =�O�a�s�ϗ��� ��������'�9�K� ]�o������������� ����+�5GYk �������� 1CUgy� ������	/# /?/Q/c/}s/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�?��?�?O/ �$E�NETMODE �1N~%��  + + �&%HOZK*@RROR�_PROG %�7J%%&�O�IxETA�BLE  7K��/�O�O_WxBSE�V_NUM FB?  �AA=P�xA_AUTO_ENB  dE?CuDw_NORQ O7K�YA<R  *�*�P��P��P��PHP�+�P�_�_�_nTFLsTRZ_lVHIS9S�)!?@g[_ALM �1P7K �&$�\% +�_no�o�o��o�o�o�__2RtP  7K�QZBz*@�TCP_VER �!7J!�O�o$E�XTLOG_RE�Qf�eY_sSI�ZhZtSTK�y��U�\rTOL � )!Dzb�{A Zt_BWD�``�p�V�q_B�sDI�qw Q~%�sxXD)!�{STEP���*@0�OP_DO��(AFDR_GR�P 1R7I�Qd �	��Z@��n&����c?���$,MT�� ��$ ���ن�������
� C�.�g�R���v���������К@م�@���?�$lA�`��
 K�&I)!�@�sW�`֟{�f�����A@/�~��@�33@�Ǡ	ˣ��@¡毄������F@ 5�E���@�5�%��L��FZ!D�`��D�� BT���@�����?� y ��#�6������5�Zf5�ES�����%9��m�*��pg����7�t��� �ۄ�KFEATURE S~%��p^AAr?cTool �)"�Englis�h Dictio�nary*�4D �Standard�#�Analog �I/O"�A5�e �Shiftw�rc� EQ Prog�ram Sele�ct��Softp�ar�ǝ�Weld���cedures<���Core���Ramping_˷uto��wa�U�pdate(�ma�tic Back�up(�V�ground Edit �~-�Camerar�=Fv�Cellr�{�nrRndIm[����ommon calib UI��F��sh������c��	���ne�	�ty���s����nt���M�onitor=�n�tr�eliab<��)�DHCP˒��ata Acqu�ish��iagn�osR�o���ocu�ment Vie�wet��ua��h�eck Safesty��-�han��o Rob��rv��q!���)�F�s��F����-�xt we�avS�ch%�xt�. DIO��nf�i"�|�end.�E�rrs�L���i�s���rm��� �p'�F�CTN Menu������TP In���fac�-�Ge�n��l��Eq L��8igE'9m��p Mask Ekxc*�gr�HT% >��xy Sv��igh-Spe.��Ski�ԍ����m�municQ�on��Hour ���s�(connX�2��ncr' str�u>��
!e���J���-�KAREL �Cmd. L� u�a�XRun-Tiq�EnvN��:�u+U�sS�S/W*�License������Book(S�ystem)'�M�ACROs,�/�OffseZ�MM�Rm�i���Mech/Stop��t����"�i���1&x.�o��S�D.od��wit���g(i���.�ƅ+O�ptm�/#��fi�l��'g��ul�ti-T  �+�O�RNTBASE �Fun+-�PCM3 f"8(�Po��� �I=Regi�r��,6ri��!9~9p��Nu����8��Ad�ju� �>���=t�atu}1�?��,�R�DM0�ot;�scgoveD�)Eea� �q�Freq An;ly��Rem' ��nR�)E5B5�9�ues�ńGo��r )�?SNPX b�#�;SN% Cli���ND��P rC��OU� 8$�P�Eo�t ssag յE���O!p1 0��V^/I&]U�MILIB�_`RP� Firm9�p^P�Accn�v�TPsTX��^Teln�`�_aQ��q]or�@ Simular���!fu��P8�XZm�t��#&��ev.]U�1�ri��_US�B po����iP��a��fR EV�NT�o�`nexcept.�j@W4�ej�P�VC��r��-(�V��.r�_?u�K9{S��@SC�UqSGE,�|uUI&�W��8�|b PlF�~5� ��� (���������6�uZDT Ap�pl�'��f�s�G�rid9AplayPm�mPZԇ�R%r.R������F� A�20�0i��c�larm Cause/h@�edE�Ascii���Load��1�U3plG���yc��~0�0�`� RAe`��<�yQ�NRTL�_4�nline Hel��-6',6{0x1���tr"�64MB �DRAM���FR!O �����c� PB� .'�mai���K��RR�6L��Sup��b�!}9à��} cr�oL4C�E��9vrt�4C&�����.�@� m�d�v�������ٿп ����3�*�<�i�`� rϟϖϨ��������� �/�&�8�e�\�nߛ� �ߤ�����������+� "�4�a�X�j���� ����������'��0� ]�T�f����������� ������#,YP b������� �(UL^� �������/ /$/Q/H/Z/�/~/�/ �/�/�/�/�/?? ? M?D?V?�?z?�?�?�? �?�?�?O
OOIO@O ROOvO�O�O�O�O�O �O___E_<_N_{_ r_�_�_�_�_�_�_o ooAo8oJowono�o �o�o�o�o�o�o =4Fsj|�� ������9�0� B�o�f�x�������ȏ ҏ�����5�,�>�k� b�t�������ğΟ�� ��1�(�:�g�^�p� ��������ʯ��� � -�$�6�c�Z�l����� ����ƿ����)� � 2�_�V�hϕόϞϸ� ��������%��.�[� R�dߑ߈ߚߴ߾��� ����!��*�W�N�`� ������������ ��&�S�J�\����� ������������ "OFX�|�� ����K BT�x���� ��///G/>/P/ }/t/�/�/�/�/�/�/ ???C?:?L?y?p? �?�?�?�?�?�?	O O O?O6OHOuOlO~O�O �O�O�O�O_�O_;_ 2_D_q_h_z_�_�_�_ �_�_o�_
o7o.o@o modovo�o�o�o�o�o �o�o3*<i` r������� �/�&�8�e�\�n��� ������ȏ�����+� "�4�a�X�j������� ��ğ����'��0� ]�T�f����������� ����#��,�Y�P� b�|����������� ���(�U�L�^�x� �ϯϦϸ�������� �$�Q�H�Z�t�~߫� �ߴ��������� � M�D�V�p�z���� �������
��I�@� R�l�v����������� ��E<Nh r������ A8Jdn� �����/�/ =/4/F/`/j/�/�/�/ �/�/�/?�/?9?0? B?\?f?�?�?�?�?�?��?�?�1  �H541�3A2�FR782 G50� EJ614DG76^ EAWSP,G1[G�RCRPH8\FTU�gFJ545DH[FV�CAM ECLIOv�FRI�GUIF,F=6�GCMSC�HgF�STYLDG2�FC�NRE,F52[FR�63+GSCH EDwOCVLVCSU E�ORSFR869�DG0OG88FEI�O�FR547FR6=9[FESET�GrG�JqIWMG�G�WM�ASK EPRXY�X7 FOC�F�P3ИH7F�PCH3fJ6�BH53{VHEhLC�H�VOPL�VJ5m0/fPS�gMCfG�`�W55OFMDS�W�g"gOP"gMP�R�F<PSh0CFOR[BS fCM�G0wl�POG50Sg51�G�51Ox0�FPRSv�W69fFRD�F�FREQ,FMCN�VmXH93CFSN�BA�GFgSHLBbVM�w<P3WNN_h�2CFHTCgFTMqIV4@{VTPA�FoTPTX(�EL�vĘ`{W86G4@FJ9�5�FTUT#g95�fUEV�VUEC��VUFR�FVCC�ψOFVIPVC;SCW�CSG'VaP�I�hOFWEBgFH�TTgG62WWIO��Ry�CG:�IG��IPGvIRCvVDG"gH75�FWR66��7�WRMz2/fR]j4f��OF��@FNVD�VD0���F�ALO�VC[TO�GNNfM}x�OLXEND,FLڇFVR�E�8���� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p�� ����� ��$� 6�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r����������̿޿���  H54�1��2#�R78�2$�50$�J61�4T�76$�AWSuP4�1s�RCRd��8t�TU��J54y5T�s�VCAM$�oCLIO��RI���UIF4�6��CM�SC4܃�STYLzT�2��CNRE4ʻ52s�R633�S{CH$�DOCV��wCSU$�ORS�ʯR869T�0c�8�8#�EIOC�R5�4C�R69s�ES�ET�˒�J��WMyG$��MASK$ɯPRXYd�7$�O	C�`�3��C�`�S�m3��J6R�53���H�LCH��OP�L��J50��PS�b�MC��p�c�55�c�MDSW����OP��MPRڠ���0S�ORBS��C�M#�0`�c�50��51��51c0n��PRSS�69���FRD��FREQ�4�MCNT���H9=3S�SNBA$��/SHLBT�M2��֓�NN#�2S�HTC��TMIc�@����TPAC�TPTXF�EL�
p���8B��@�#�J95��TU�T��95��UEV�S�UEC��UFR���VCCc,O��V�IPc�CSC�C�SG����Id�c�W�EB��HTT��6���WIO�*R�C�G�+IG�+IPGn#
IRCc�DG��wH75��R66�;U7B�Ra2��R!��4��0c�0�#�NV�DS�D0�;F!LA�LO��CTO��N�N��M�OLR�E�ND4�Lr+FVR C�ȺO�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p�����@����ʿܿ� ���STD�LANG(�#�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K]�o��RBT'�OPTN�����
+DPN&�"/4/F/X/j/|/���/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?� ?2?D?V?h?z?  ��?�?�?�?�?�?�=�99E�$FE�AT_ADD ?_	���/A7@?  	�8@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r����������� ��&�8�J�\�n��� ���������������""DDEMO �S/I    �8i_q���� ��
-7d [m������ /�/)/3/`/W/i/ �/�/�/�/�/�/?�/ ?%?/?\?S?e?�?�? �?�?�?�?�?�?O!O +OXOOOaO�O�O�O�O �O�O�O�O__'_T_ K_]_�_�_�_�_�_�_ �_�_�_o#oPoGoYo �o}o�o�o�o�o�o�o �oLCU�y �������� �H�?�Q�~�u����� ���������D� ;�M�z�q��������� �ݟ�	��@�7�I� v�m���������ٯ ���<�3�E�r�i� {�������޿տ�� �8�/�A�n�e�wϤ� �ϭ����������4� +�=�j�a�sߠߗߩ� ���������0�'�9� f�]�o�������� ������,�#�5�b�Y� k��������������� ��(1^Ug� �������$ -ZQc��� ����� //)/ V/M/_/�/�/�/�/�/ �/�/�/??%?R?I? [?�??�?�?�?�?�? �?OO!ONOEOWO�O {O�O�O�O�O�O�O_ __J_A_S_�_w_�_ �_�_�_�_�_ooo Fo=oOo|oso�o�o�o �o�o�oB9 Kxo����� ����>�5�G�t� k�}�������͏׏� ���:�1�C�p�g�y� ������ɟӟ ���	� 6�-�?�l�c�u����� ��ůϯ����2�)� ;�h�_�q��������� ˿����.�%�7�d� [�mϚϑϣϽ����� ����*�!�3�`�W�i� �ߍߟ߹��������� &��/�\�S�e��� ����������"�� +�X�O�a��������� ��������'T K]������ ��#PGY �}������ ///L/C/U/�/y/ �/�/�/�/�/�/?	? ?H???Q?~?u?�?�? �?�?�?�?OOODO ;OMOzOqO�O�O�O�O �O�O
___@_7_I_ v_m__�_�_�_�_�_ o�_o<o3oEoroio {o�o�o�o�o�o�o 8/Anew� �������4� +�=�j�a�s�����ď ��͏����0�'�9� f�]�o���������ɟ �����,�#�5�b�Y� k���������ů�� ��(��1�^�U�g��� ������������$� �-�Z�Q�c�}χϴ� �Ͻ������� ��)� V�M�_�y߃߰ߧ߹� ��������%�R�I� [�u��������� ����!�N�E�W�q� {������������� JASmw� ����� F=Ois��� ���///B/9/ K/e/o/�/�/�/�/�/ �/?�/?>?5?G?a? k?�?�?�?�?�?�?O �?O:O1OCO]OgO�O �O�O�O�O�O _�O	_ 6_-_?_Y_c_�_�_�_ �_�_�_�_�_o2o)o ;oUo_o�o�o�o�o�o �o�o�o.%7Q [���������*�!�M�  D�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� 1CUgy� ������	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? m??�?�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_ �_�_�_�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K ]o������ ���#�5�G�Y�k� }�������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w��� �����������+� =�O�a�s��������� ������'9K	  LQg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� ����#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{�������������@��/APU Hk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����������/�A�S���$FEAT_DEMOIN  X������X�k�I�NDEXx�����k�ILECOMP T��������f���SETUP2 U���Â�  N� �_AP2B�CK 1V�� � �)T�"�1�%�U�X���C���V� ���;�П_�ݟ��� *���N�`����� ��I�ޯm�����8� ǯ\��i���!���E� ڿ�{�ϟ�4�F�տ j����Ϡ�/���S��� w���߭�B���f�x� ߜ�+�����a��߅� �,��P���t��� ��9���]������(� ��L�^��������� G���k� ��6�� Z��~��C� �y�2D�h ����Q�u 
//�@/�d/v// �/)/�/�/_/�/�/?��/%?N?ȉ��P �� 2�*.VRU?�?0*�?�?
30�?�?�%�0PC�?#O>0FR6:OON�?sOKT���O�O�8E�O�Lz�dO�O�&G*.F�?*_1	:C�_W\�O{_
[ST�M�_�_7B=@�_�]j_�_
[H�_2o�W op�_�_�oZGIF�o��o�U�oaosoZJPG<�U(�o�o��JJS��0�Rs�j%
JavaScript�CS�C��V0��� %Casca�ding Sty�le Sheet�so�� 
ARGN?AME.DT��<�P\��p��q������DISP*��.ބ9���	�i��w�#�
TPEIN�S.XML��Ώ:�\��x�ځCust�om Toolb�ar��*�PASS�WORDn��.F�RS:\>���_�P�assword ?Config��/ ȯW�����4?"���F� X��|������A�ֿ e�������0Ͽ�T�� Mϊ�Ϯ�=�����s� ߗ�,�>���b��φ� �'߼�K���o���� ��:���^�p��ߔ�#� ����Y���}����� H���l���e���1��� U������� ��DV ��z	�-?�c ���.�R�v ��;��q/ �*/��`/��// }/�/I/�/m/??�/ 8?�/\?n?�/�?!?�? E?W?�?{?O�?	OFO �?jO�?�O�O/O�OSO �O�O�O_�OB_�O�O x__�_+_�_�_a_�_ �_o,o�_Po�_to�o o�o9o�o]ooo�o (�o!^�o�� �G�k ���6� �Z��������C� ���y����2�D�ӏ h�������-�Q�� u������@�ϟ9�v� ���)���Я_����� �*���N�ݯr��� ��7�̿[�ſϑ�&� ��J�\�뿀�Ϥ϶� E���i��ύϟ�4����$FILE_D�GBCK 1V���!���� < �)
�SUMMARY.�DG>���MD:�r߲���Dia�g Summar�y����
CONSLOG�ߋߝ���6����Consol�e log7��	?TPACCN,���%y����TP �Accounti�nX���FR6:�IPKDMP.ZIP����
�;������Excepti�on?����MEMCHECK�������J�Memor?y Data����3l�)	FTAP)�����L��mment TB�DG�L >I)�ETHERNE�T<�΁�����Ethernet� N�figura�^���1DCSVR�F;!3L��%� verif�y allO�M�.cDIFF�D*<���%fdiff����>CHG01����V/a�~/�- )2L/3/E/�/�{/��/"3�/�/�/^?� �/�?6VT�RNDIAG.LAS�?;?M?�?���1� Ope� Lo�g ��nosti�c��:�)VwDEV�2DAT�?��?�?�?bVis~ADeviceOKIMG�21�AOSO��O�#~DImag܊OKUP/@ES�.O�OFRS:\�._o]��Upda�tes List�o_���@FLEXEVEN��O�O�_�a�Q UIF �Evb	@�_  ,��t)
PSRBWLD.CMo���ZR6oq_K�PS�_ROBOWEL|h�:GIGE	�Oo�_�o��Gig�EXo�N�A��)�aHADOW��o�o�o|��Sh�adow Cha�nges��a��<rRCMERR�tYk ����pC�FG Errorބ@tail� M�A����pSGLIB�����rI�� St� A-�>�7�)r�ZD�o���o����ZD@a�d��3� <rNO�TI�������Notific�3�(f�AG����� ���;���_�� ��$���H�ݯ�~�� ��7�I�دm����� � ��ǿV��z��!ϰ� E�Կi�{�
ϟ�.��� ��d��ψ�߬�*�S� ��w�ߛ߭�<���`� ����+��O�a��� ����8����n�� ��'�9���]������ "���F�����|��� 5��Bk���� �T�x�C �gy�,�P ���/�?/Q/� u//�/�/:/�/^/�/ ?�/)?�/M?�/Z?�? ?�?6?�?�?l?O�? %O7O�?[O�?O�O O �ODO�OhO�O_�O3_ �OW_i_�O�__�_�_ R_�_v_oo�_Ao�_ eo�_ro�o*o�oNo�o �o�o�o=O�os ��8�\�� �'��K��o���� ��4�ɏۏj�����#� 5�ďY��}������ B�ןf������1��� U�g����������P� �t�	����?�ίc� 򯇿��(���L������Ϧ�;�M��$F�ILE_FRSP�RT  ���1�����\�MDONLY �1Vp�(� 
� �)MD:_�VDAEXTP.�ZZZN��������6%NO B�ack filey ��(�S�6)ܿ 7���[�$�hߑ�ֿ�� D�����z���3�E� ��i��ߍ��.���R� ��v������A���e� w����*�����`��� ��+��O��s ��8�\�� '�K]�����`�VISBCK���x���*.VD��/pFR:\��ION\DAT�A\��pV�ision VD �./<v/�/��/� �/_/�/?�/*?�/N? `?�/�??�?7?I?�? m?OO�?8O�?\O�? mO�O!O�OEO�O�O{O _�O4_�O�Oj_�O�_ �_[_�_S_�_w_�_o �_Bo�_foxoo�o+o��oOoao�oV�LUI�_CONFIG �Wp��{O $ �c��{p� Xj|����y@p|x�o��� �2� B��e�w�������D� �������+�O� a�s�������@�͟ߟ ���'���K�]�o� ������<�ɯۯ��� �#���G�Y�k�}��� ��8�ſ׿����� ��C�U�g�yϋϝ�4� ��������	ߠ��?� Q�c�u߇�߽߫��� ������)�;�M�_� q����������� ���%�7�I�[�m�� ��������������� !3EWi{� ������/ ASe�v��� ��z//+/=/O/ a/��/�/�/�/�/�/ v/??'?9?K?]?�/ �?�?�?�?�?�?r?�? O#O5OGOYO�?}O�O �O�O�O�OnO�O__ 1_C_U_�Oy_�_�_�_ �_X_�_�_	oo-o?o �_couo�o�o�o�oTo �o�o);�o_ q����P�� ��%�7��[�m�� ������L�ُ���� !�3�ƏW�i�{��������A�͐x��ʓ��$FLUI_DA�TA X��}���D���RESULT �2Y��#� ��T�/wiz�ard/guid�ed/steps/Expertٟ Z�l�~�������Ưد�������Co�ntinue w�ith G7�ance�W�i�{��������ÿտ����� �˒-̑��<�0 �M�<�����\��.�psϧϹ� ��������%�7�I� [�m�,�M��ߦ߸��� ���� ��$�6�H�Z�@l�~�\�N�`�r���torch����� �*�<�N�`�r����� ����y�����& 8J\n��������������wproc��HZl~ �������/ ��2/D/V/h/z/�/�/ �/�/�/�/�/
??���7?{���@�T�imeUS/DST&?�?�?�?�?�?O�O,O>OPObO%�EnablE��O�O�O �O�O�O__&_8_J_\_n_˒8�F?�_j?|?�624�?�_o "o4oFoXojo|o�o�o �oqO�O�o�o0 BTfx�����_�_�_�_w�-�?�Region�R�d� v���������Џ����!�America<@�R�d�v��� ������П����!��qy��P��$��2Edi�������ʯ ܯ� ��$�6�H�Z��+ Touch �Panel �� �(recommen��)h�����ѿ� ����+�=�O�a� ���0�B���f�x��2acces/����� /�A�S�e�w߉ߛ߭��,Connec�t to Network������ )�;�M�_�q������$���p�ϚϬ���\!�ϐ0Introduct>�Q�c� u���������������  /);M_q� ������ 0?��0
��R# �������/ /(/:/L/^/�/�/ �/�/�/�/�/ ??$?6?H?Z?�x3P:H�?l�?�?�?O O+O=OOOaOsO�O�O �Oh/�O�O�O__'_ 9_K_]_o_�_�_�_�_ v?�?�?�_�?#o5oGo Yoko}o�o�o�o�o�o �o�o�O1CUg y������� 	��_*��_N�ou��� ������Ϗ���� )�;�M�_�p������� ��˟ݟ���%�7� I�[��|�>���b�ǯ ٯ����!�3�E�W� i�{�������p�տ� ����/�A�S�e�w� �ϛϭ�l��ϐ��ϴ� ��+�=�O�a�s߅ߗ� �߻��������¿'� 9�K�]�o����� ��������� ���D� V��}����������� ����1CU� y������� 	-?Q�Z�4� ~�j����// )/;/M/_/q/�/�/�/ f�/�/�/??%?7? I?[?m??�?�?b� ��?�?�!O3OEOWO iO{O�O�O�O�O�O�O �O�/_/_A_S_e_w_ �_�_�_�_�_�_�_�? �?�?�?LoOso�o�o �o�o�o�o�o' 9K
_o���� �����#�5�G� Y�o*o<o��`oŏ׏ �����1�C�U�g� y�����\��ӟ��� 	��-�?�Q�c�u��� ����j�|���𯲏� )�;�M�_�q������� ��˿ݿ￮� �%�7� I�[�m�ϑϣϵ��� �����ϼ���B�� i�{ߍߟ߱������� ����/�A�S�d�w� ������������ �+�=�O��p�2ߔ� V߻�������' 9K]o���d� ����#5G Yk}��`���� ����/1/C/U/g/ y/�/�/�/�/�/�/�/ �?-???Q?c?u?�? �?�?�?�?�?�?�O �8OJO?qO�O�O�O �O�O�O�O__%_7_ I_?m__�_�_�_�_ �_�_�_o!o3oEoO NO(Oro�o^O�o�o�o �o/ASew ��Z_����� �+�=�O�a�s����� Vo�ozoďo�'� 9�K�]�o��������� ɟ۟ퟬ�#�5�G� Y�k�}�������ůׯ 鯨���̏ޏ@��g� y���������ӿ��� 	��-�?���c�uχ� �ϫϽ��������� )�;�M���0���T� ����������%�7� I�[�m���Pϵ��� �������!�3�E�W� i�{�����^�p߂��� ��/ASew ��������� +=Oas�� �������/�� 6/��]/o/�/�/�/�/ �/�/�/�/?#?5?G? X/k?}?�?�?�?�?�? �?�?OO1OCO/dO &/�OJ/�O�O�O�O�O 	__-_?_Q_c_u_�_ �_X?�_�_�_�_oo )o;oMo_oqo�o�oTO �oxO�o�O�o%7 I[m���� ���_�!�3�E�W� i�{�������ÏՏ� �o��o,�>��e�w� ��������џ���� �+�=��a�s����� ����ͯ߯���'� 9���B��f���R��� ɿۿ����#�5�G� Y�k�}Ϗ�N������� ������1�C�U�g� yߋ�J���n����ߤ� 	��-�?�Q�c�u�� ����������� )�;�M�_�q������� �������߮�����4 ��[m���� ���!3��W i{������ �////A/ $ �/H�/�/�/�/�/? ?+?=?O?a?s?�?D �?�?�?�?�?OO'O 9OKO]OoO�O�OR/d/ v/�O�/�O_#_5_G_ Y_k_}_�_�_�_�_�_ �?�_oo1oCoUogo yo�o�o�o�o�o�o�O �O*�OQcu� �������� )�;�L_�q������� ��ˏݏ���%�7� �oX�|�>����ǟ ٟ����!�3�E�W� i�{���L���ïկ� ����/�A�S�e�w� ��H���l�ο����� �+�=�O�a�sυϗ� �ϻ����Ϟ���'� 9�K�]�o߁ߓߥ߷� ���ߚ��߾� �2��� Y�k�}�������� ������1���U�g� y��������������� 	-��6��Z� F����� );M_q�B�� ����//%/7/ I/[/m//>�b�/ �/��/?!?3?E?W? i?{?�?�?�?�?�?� �?OO/OAOSOeOwO �O�O�O�O�O�/�/�/ �/(_�/O_a_s_�_�_ �_�_�_�_�_oo'o �?Ko]ooo�o�o�o�o �o�o�o�o#5�O __z<_���� ����1�C�U�g� y�8o������ӏ��� 	��-�?�Q�c�u��� FXj̟���� )�;�M�_�q������� ��˯��ܯ��%�7� I�[�m��������ǿ ٿ���������E�W� i�{ύϟϱ������� ����/�@�S�e�w� �ߛ߭߿�������� �+��L��p�2ϗ� �����������'� 9�K�]�o���@ߥ��� ��������#5G Yk}<�`���� ��1CUg y�������� 	//-/?/Q/c/u/�/ �/�/�/�/��/�? &?�M?_?q?�?�?�? �?�?�?�?OO%O� IO[OmOO�O�O�O�O �O�O�O_!_�/*?? N_x_:?�_�_�_�_�_ �_oo/oAoSoeowo 6O�o�o�o�o�o�o +=Oas2_|_ V_���_���'� 9�K�]�o��������� ɏ�o����#�5�G� Y�k�}�������ş� �����C�U�g� y���������ӯ��� 	��ڏ?�Q�c�u��� ������Ͽ���� )�����n�0��ϧ� ����������%�7� I�[�m�,��ߣߵ��� �������!�3�E�W� i�{�:�L�^������ ����/�A�S�e�w� ��������~����� +=Oas�� ���������� 9K]o���� ����/#/4G/ Y/k/}/�/�/�/�/�/ �/�/??�@?d? &�?�?�?�?�?�?�? 	OO-O?OQOcOuO4/ �O�O�O�O�O�O__ )_;_M___q_0?�_T? �_x?z_�_oo%o7o Io[omoo�o�o�o�o �O�o�o!3EW i{�����_� �_���oA�S�e�w� ��������я���� ��o=�O�a�s����� ����͟ߟ���� ��B�l�.������� ɯۯ����#�5�G� Y�k�*�������ſ׿ �����1�C�U�g� &�p�J��Ͼπ����� 	��-�?�Q�c�u߇� �߽߫�|������� )�;�M�_�q���� ��xϊϜϮ����7� I�[�m���������� ��������3EW i{������ ����� �b$� �������/ /+/=/O/a/ �/�/ �/�/�/�/�/??'? 9?K?]?o?.@R�? v�?�?�?O#O5OGO YOkO}O�O�O�Or/�O �O�O__1_C_U_g_ y_�_�_�_�_�?�_�? o�?-o?oQocouo�o �o�o�o�o�o�o (o;M_q��� �������_4� �_X�o�������Ǐ ُ����!�3�E�W� i�(������ß՟� ����/�A�S�e�$� ��H���l�n����� �+�=�O�a�s����� ����z�߿���'� 9�K�]�oρϓϥϷ� v��Ϛ����ҿ5�G� Y�k�}ߏߡ߳����� �����̿1�C�U�g� y������������ 	������6�`�"߇� ������������ );M_��� ����%7 I[�d�>���t� ���/!/3/E/W/ i/{/�/�/�/p�/�/ �/??/?A?S?e?w? �?�?�?l~��O �+O=OOOaOsO�O�O �O�O�O�O�O_�/'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o�?�?�? VoO}o�o�o�o�o�o �o�o1CU_ y������� 	��-�?�Q�c�"o4o Fo��joϏ���� )�;�M�_�q������� f��ݟ���%�7� I�[�m��������t� ֯������!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� Ư(��L��s߅ߗ� �߻���������'� 9�K�]�ρ���� ���������#�5�G� Y��z�<ߞ�`�b��� ����1CUg y���n���� 	-?Qcu� ��j�����/� )/;/M/_/q/�/�/�/ �/�/�/�/?�%?7? I?[?m??�?�?�?�? �?�?�?�/�*OTO /{O�O�O�O�O�O�O �O__/_A_S_?w_ �_�_�_�_�_�_�_o o+o=oOoOXO2O|o �ohO�o�o�o' 9K]o���d_ �����#�5�G� Y�k�}�����`oro�o �o���o�1�C�U�g� y���������ӟ��� ��-�?�Q�c�u��� ������ϯ���ď ֏�J��q������� ��˿ݿ���%�7� I��m�ϑϣϵ��� �������!�3�E�W� �(�:���^������� ����/�A�S�e�w� ���ZϬ�������� �+�=�O�a�s����� ��h���������' 9K]o���� ����#5G Yk}����� ����/��@/g/ y/�/�/�/�/�/�/�/ 	??-???Q?u?�? �?�?�?�?�?�?OO )O;OMO/nO0/�OT/ VO�O�O�O__%_7_ I_[_m__�_�_b?�_ �_�_�_o!o3oEoWo io{o�o�o^O�o�O�o �o�_/ASew ��������_ �+�=�O�a�s����� ����͏ߏ�o�o�o �H�
o��������� ɟ۟����#�5�G� �k�}�������ůׯ �����1�C��L� &�p���\���ӿ��� 	��-�?�Q�c�uχ� ��X����������� )�;�M�_�q߃ߕ�T� f�x����߮��%�7� I�[�m������� ������!�3�E�W� i�{������������� ��������> �ew ������� +=��as�� �����//'/ 9/K/
.�/R�/ �/�/�/�/?#?5?G? Y?k?}?�?N�?�?�? �?�?OO1OCOUOgO yO�O�O\/�O�/�O�/ 	__-_?_Q_c_u_�_ �_�_�_�_�_�__o )o;oMo_oqo�o�o�o �o�o�o�o�O�O4 �O[m���� ����!�3�E�o i�{�������ÏՏ� ����/�A� b�$ ��HJ���џ���� �+�=�O�a�s����� V���ͯ߯���'� 9�K�]�o�����R��� v�ؿ꿮��#�5�G� Y�k�}Ϗϡϳ����� �Ϩ���1�C�U�g� yߋߝ߯������ߤ� �ȿ�<���c�u�� ������������ )�;���_�q������� ��������%7 ��@��d�P�� ���!3EW i{�L����� �////A/S/e/w/ �/HZl~�/�? ?+?=?O?a?s?�?�? �?�?�?�?�OO'O 9OKO]OoO�O�O�O�O �O�O�O�/�/�/2_�/ Y_k_}_�_�_�_�_�_ �_�_oo1o�?Uogo yo�o�o�o�o�o�o�o 	-?�O_"_� F_������� )�;�M�_�q���Bo�� ��ˏݏ���%�7� I�[�m����P��t ֟����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ㿢�� Ɵ(��O�a�sυϗ� �ϻ���������'� 9���]�o߁ߓߥ߷� ���������#�5��� V��z�<�>������ ������1�C�U�g� y���J߯��������� 	-?Qcu� F�j����� );M_q��� �����//%/7/ I/[/m//�/�/�/�/ �/���?0?�W? i?{?�?�?�?�?�?�? �?OO/O�SOeOwO �O�O�O�O�O�O�O_ _+_�/4??X_�_D? �_�_�_�_�_oo'o 9oKo]ooo�o@O�o�o �o�o�o�o#5G Yk}<_N_`_r_� �_���1�C�U�g� y���������ӏ�o�� 	��-�?�Q�c�u��� ������ϟ០�� &��M�_�q������� ��˯ݯ���%�� I�[�m��������ǿ ٿ����!�3��� �x�:��ϱ������� ����/�A�S�e�w� 6��߭߿�������� �+�=�O�a�s��D� ��h��������'� 9�K�]�o��������� ��������#5G Yk}����� �������CUg y������� 	//-/��Q/c/u/�/ �/�/�/�/�/�/?? )?�J?n?02?�? �?�?�?�?OO%O7O IO[OmOO>/�O�O�O �O�O�O_!_3_E_W_ i_{_:?�_^?�_�_�O �_oo/oAoSoeowo �o�o�o�o�o�O�o +=Oas�� ����_�_�_�$� �_K�]�o��������� ɏۏ����#��oG� Y�k�}�������şן ������(��L� v�8�������ӯ��� 	��-�?�Q�c�u�4� ������Ͽ���� )�;�M�_�q�0�B�T� f��ϊ�����%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{��������� �ϸ����A�S�e�w� �������������� ��=Oas�� �����' ����
�l.���� ����/#/5/G/ Y/k/*|/�/�/�/�/ �/�/??1?C?U?g? y?8�?\�?��?�? 	OO-O?OQOcOuO�O �O�O�O�O�?�O__ )_;_M___q_�_�_�_ �_�_�?�_�?o�?7o Io[omoo�o�o�o�o �o�o�o!�OEW i{������ ����_>� ob�$o &�������я���� �+�=�O�a�s�2�� ����͟ߟ���'� 9�K�]�o�.���R��� Ư������#�5�G� Y�k�}�������ſ�� �����1�C�U�g� yϋϝϯ��π�ʯ�� ���گ?�Q�c�u߇� �߽߫��������� ֿ;�M�_�q���� ������������� ��@�j�,ߑ������� ������!3EW i(������ �/ASe$� 6�H�Z��~���/ /+/=/O/a/s/�/�/ �/�/z�/�/??'? 9?K?]?o?�?�?�?�?��?���OE�$�FMR2_GRP� 1ZE�� �C4 w B�� 	 � �VOhLS@F@ ~EE���B~A�:{A��L�FZ!D��`�D�� BT��@��ÖM�?�  �O�<S@6�����B��5�Zf5�ESQ��MA�  _0[B�HT�@JQ@�33K@�TPXS�<RDx_�]S@@OQ�_�N�_��_RA<�z�<��ڔ=7�<��
;;�*�<����M8ۧ�9�k'V8��8����7ג	8(���_?o�_<ouo�`o�o�o�o�',B_C_FG [9KThB��o/�iNO {9J
F0cq� hp�lRM_CHKTYP  )A�� A@C@�0+AROM�~p_MIN�p�#����p�oPX,@S�SB�c\E TF��%�s����eTP_DEF_OW  �$�AC$�IRCOM��p5��$GENO�VRD_DO�v��!b�THR�v dz�dh�_ENBT�{ h�RAVC2Cu]�w�p �vE � ��o$��L2�C�nfZ �ȁOU5@c9LkqfH9�fE<�p�O��d����ԟ��#C�  D +�1���L�\�@OAC�B�gAI�iI���ɀSMT2Cd։E@�p�'��$HOSTC��b1e9I�p�\�/R@ MC�$?�����&  2�7.0M�16�  e-�z��������� h�����:�ѿ˳�	anonymous>�l�~ϐϢϴ��"��Q@����+�-� �a�B�T�f�xߊ�Ϳ ��������ߡ�K�,� >�P�b�t�������� �����5��(�:�L� �	������������� � $6H���� ����������  c�DVhz� ��������
// _q���m/��/ �/�/�/�/7?*?<? N?`?�/���?�?�? �?�?3/E/W/i/k?\O �/�O�O�O�O�O?�O �O_"_4_WO�?N_|_ �_�_�_�_OO+O�_ ?_0osOTofoxo�o�o �O�o�o�o�oo]_ >Pbt���_�_ �_��Go(�:�L� ^��o��������ʏ� o�1�$�6�H�Z���~ߡENT 1f�?�  P!鏫�  ����֟ş ������B��N�)� w���_�����䯧�� ˯,���b�%���I� ��m�ο�����ǿ(� �L��p�3�iϦϕ� �ύ��ϱ������� G�l�/ߐ�Sߴ�w��� ���߿���2���V���z�=�QUICCA0��c�u����1������&���2'����v�!ROUTE�Rw�S�e���!P�CJOG����!�192.168�.0.10���C�AMPRT��!�1 >%RT��BT� !S�oftware �Operator? Panel��{�NAME �!��!ROBO�0S_CFG �1e�� ��Auto-s�tarted�tFTP���ޏ ����/#/5/~� Y/k/}/�/��/F/�/ �/�/??1?�pw� �|?�/��?�?�?�? �?�/O0OBOTOfO�? O�O�O�O�O�O�O� ���qOG_�?�_�_ �_�_�_�O�_oo(o :o]_�_po�o�o�o�o �o__1_C_Eo6y_ Zl~��eo�� ���1�D�V�h� z������o�o��� 
�M.�@�R�d�v�9� ������П������ *�<�N�`�r���Ǐُ ���ޯ!���&�8� ��\�n�������ǯI� ÿ����"�4�w��� ��������������� ���Ͽ0�B�T�f�x� ��߮���������� K�]�oρσ�t�Ϙ� ����������(� :�L�o���������������_ERR �g&����PDU�SIZ  q�^ڏ��>$WR�D ?eR�� � guestq�dv�����SCD_GR�OUP 3he ui{�IFTw$PAOMPw _SH�EDS $CC�OM��TTP_A�UTH 1i� <!iPen�dan���q��n1!KAREL�:*���KC�//'/�VISION SET� �/\/m6!�/�/�/� �/�/�/�/7?? ?m?�D?V>�CTRL Kj�8q�
q��FFF9E3�y?P�FRS:D�EFAULT�<�FANUC W�eb Server�:�2R�L^�<�YOkO}O�O�O�O��W�R_CONFIGw k�?��?��IDL_C_PU_PC@q�sB�S�%P BHU�MIN\�)UGNR_IO��2q�	�PNPT_SIM�_DO[Ve[STAL_SCRN[V� ��6oQTPMODNTOL�We[>ARTY|X%QjVy ��ENB�W�
SO�LNK 1l  -o?oQocouo�o�o�bMASTEZP�ijUOSLAVE� m�eRAM�CACHE�o�RO>�O_CFG�oc�sUO� rCMT_OP@]R
Os�YCL�o+u�0_A�SG 1n�G>
 �o����� �*�<�N�`�r���������k�rNUM1�	
rIP�owR?TRY_CNZ+u��Q_UPD1,a�b r8pro�n�� g�� PRCA_�ACC 2p��  Wi! ;^kq�6���1�q�5�3 R�૟���3̜}�BUF�001 2q�=� h/u0  �u0h@�O�`��o���������������Z���i~�~��!~�-[,`[d���e	����)���8��I��X��i���x���������������ʦ�٦��Z����f&�&�U+&�:&�L&�[&�Ul&�{&��&��&�U�&��&��&��&���&���g�����.��=��N��]ꦴn��}� 8.S�8h� ���2���$�)�-�)� 5�)�=�)�E�)�M�)� U�)�]�)�e�)�m�)� u�)�}�����������������i`Ь�����½���Š ��͠��ՠ��ݠ���W�p졹����� ������������� ���%��,�1�5�1� =�1�E�1�M�1�U�1� ]�1�e�1�m�1�u�1� }�1҅�1ҍ�1ҕ�1� ��1ҥ�����ҵ��� ����Ű��Ͱ��հ�� ݰ���)�����)������3��+�2� -�;�2�=�K�2�M�[� 2�]�k�2�m�{�2�}� �Ò⍢�Ò❢��v� ����v���v�͢�� v�ݢ��v����v��� �v���v��+�q� ,�;�:�=�K�:�M�[� :�]�k�:�m�{�:�}� ��:򍲛�:򝲫�\ ���Ӻ��Ӻ�Ͳ�� ��ݲ��2����2������q2r� 4��<�5\\<\pPS]R}�HIS��t� ܛ� �2023-08-k16\+g7\A;�����Zh\�:��� 2DSW����7���������R	AS �	A��P/#/|= 3,k�}j/|/�/�/�/ �/�/�/�/?C/U/B? T?f?x?�?�?�?�?�? �??-?O,O>OPObO tO�O�O�O�O�?O�O __(_:_L_^_p_�_ �_�O�O�O�_�_ oo $o6oHoZolo��k� w�w� d{o�o(�o�9: c��cK]o]ox�������Sd  �b	 !��G��_�_ �������ŏ׏��� ��1�h�z�g�y��� ������ӟ���	�@� R�?�Q�c�u������� ��ϯ��*��)�;� M�_�q���������� ����%�7�I�[� m�ϑ�o�e��o�o �� C	��)�;� C��k�}ߏ�}� ������������ "��	 Z�g�y�׿� ����������	��-� ?�Q����������� ������)`�r� _q������ �8J\I[m ������" 4!/3/E/W/i/{/�/�/�/�/�eI_CF�G 2u�� H�
Cycle �Time�Bu{sy�Idl2��min�+R��Up�&�R�ead7DoYw+8'? ;2�#�Count�	N'um �"����<��1�aPROG��"v����� �?�?O!O3OEOWO29��eSDT_ISO�LC  ��� ��@�.J23_D�SP_ENB  ��KPЫ@INC �w�M�Ә@A  � ?�=���<�#�
�A�I:�o �A_(_��_P_��G�0GROUP �1x�K!�<A �C��_X_?��?�_��Q�_o!o�3o�_Woio{o�o��@_b[IN_AUT�O  ���J�@POSREC�C�b71��hKANJI_M�ASK�f�jKAR�ELMON y�˰?��yRok}�����.)r�3z�7��C���u�ouCL;_L�`NUM�@
���@KEYLOGG'ING�`����Q�E��0LANGUAG�E ��q���DEFAUL�T ���LG�!Y{�:72��x�@߰  8P�H [ ���'0����囿�cOU�;���
�(UT1:\�� ��.� @�W�d�v�����������(Z���LN_DISP |�O�48�_�_!�OCTOL`���Dz�0�A�A�v�GBOOK }��dޔR��ᑮ�Xٌү������,�<���P�N�*�	 ��ۉ�QmK��aO�A���_BUFF 2~N�K ���235 ݿ��R���17�'�T� K�]ϊρϓ��Ϸ��� �������#�P�G�Y�����C��DCS ��9�B�AK�����%��� ��$��IO ;2��� !Z��Q�]�m���� �����������!�5� E�W�i�}����������������8�ER_ITM�Nd�ofx ������� ,>Pbt�����p�;SEVt�`�M7TYP�N�U6/H/Z/��aR�ST(���SCRN�_FL 2�F��0����/�/�/??(?:?k/TP>��O%"}M=NGNAM�D�ǥq���UPS)�G�I� 	��E�1_�LOADPROG� %g:%	T_ARCWELDG?��MAXUALR�M%��a���E
�B�1_PR�4�` h��L�@C,�����hO���%��ODoPP �2��� �ؖ	 %/�O�O�O�O_-__ Q_<_u_X_j_�_�_�_ �_�_o�_)ooMo0o Bo�ono�o�o�o�o�o �o%[F j������� �3��W�B�{���p� ����Տ��ʏ���/� �S�e�H���t����� ���Ο��+�=� � a�L���h�z�����߯ ʯ����9�$�]�H�DBGDEF �YE��eOu�_LDXDISA�0f;6�MEMO_AP�0�E ?g;
 ��F������/��A�S�e�@FRQ_�CFG �YG6��A F�@���H�<��d%h���yϋ���B�YKL��*�/� **:(�H��-���H� S�eߒ߉ߛ��߿��� ��J�YE'� �N�<�R�`�,(�ߥ��� ��������*��N� 5�r���k������������JISC 1�g9� �P�JL� ��`K���� �_MSTR ����SCD 1�ֽ��/�S>w b������� //=/(/M/s/^/�/ �/�/�/�/�/?�/ ? 9?$?]?H?�?l?�?�? �?�?�?�?�?#OOGO 2OkOVOhO�O�O�O�O �O�O_�O_C_._g_ R_�_v_�_�_�_�_�_ 	o�_-ooQo<ouo`o �o�o�o�o�o�o�ox;�MJPT��1��i�{�w^s�MIR 1���^�p ��Lx��.s< ���?O�.q?y�3\�N�� � ���P����.��©� &��5C��o.q ���~�+yH��@�b� ��v���Ə珺�� ��ҏD�b�4�^���b� ����П��؟�+y�� ��L�^�����g�q� ��ͯk�ů����� K�-�~�����5�W�ɿ ����׿ϯ��G�-� ?�a�c�q�����g�y� �������U�;�]� ��qߓ��ߣϵ��� �߽�?���3�=��a� ������������ J�\������e�w�� ��i���������I +�|��3U��� ���E+=�_�o^pKdq��j{  �\rLT�ARM_��ju�p�xtop/$^p�METPU  �.r���]qND�SP_ADCOLx3%�>.CMNTT/ G%FNp t/E'�FSTLI�/�'MST ���/xs�� ?
4G%POSC�F�'.PRPMls/9STR 1�j}=4�q<#�
�16q �5�?�7�?�?�?�?�? �?�?.OO"OdOFOXO �O|O�O�O�O�O_�A�G!SING_CH�K  �/$MOWDAQ��jy���@UDEV 	�jz	MC:t\HOSIZE3 ��@UTASK %jz�%$123456�789 �_�U>WT�RIfp�j{ lju%�8oh+oloOm��t�SYP�Q{uVT�?SEM_INF �1��XQ`)�AT&FV0E�0uo�m)�aE0�V1&A3&B1�&D2&S0&C�1S0=�m)A#TZ�o@'tHDl�a`o�#xA������ �oC��o ,��P���� ����֏?�Q�8�u� (�:���^�p������ ��)�`�M�����>� ����˯ݯ�����Ɵ ؟�[��������� h�ٿ�������3�� ��i��.�@�����v� ������пA���e� L߉ߛ�NϿ�rτϖ� �����=�O��s�&߀��R�������m_N�ITOR� G ?��[   	EOXEC1�"3�2:�3:�4:�5:�`<�U7:�8:�9:�5� �ҟ�9��E��Q�� ]��i��u����P������2��2��U2��2��2��2��U2��2��22�3��3��3E�@QR�_GRP_SV �1��k (�A@��?������I�?�Bc��� �����Q_D��^�IO/N_DBJP�N]�!_  �� McXX?)0J�� 
cX���N _\?(cY-ud1�U�����aPL_NAME� !e��!�Default� Persona�lity (fr?om FD)G �RR2� 1�L�XL�x�hP d�"J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�2F/�? OO%O7OIO[OmOO�O�<�?�O�O�O�O __'_9_K_]_o_�_$��F�O�^
�_�_�P�_oo/oAoSo eowo�o�o�o�o�o�o �o�_�_Oas �������� �'�9�K�]�,>�� ����ɏۏ����#� 5�G�Y�k�}�������� H�6 H?�b H\��� �  ����d ܓĐ�#��E�S�Ő ���=����������� ��ٯϯ�� ��5�W�� z������	`ï��Ͽ|ῠ�:�oA���,π AH� Lɨ�'tw.������e�~� �G�� hȟ���ϰ���������
�C��R� 1��u��@ �� ����� �@D�  ��?�ěӁ�?��тA�?�6Ez  �ј���;�	l��	 ��@�? 0vw��� ���� � �� ��� J���K ��J�˷�J� �J�4�JR�<(��7'��d���S��@�;fA6�A��A1U�A��X@�O��=��N��f������T;f���X���E���*  ��  ß5��>������ҘM�?��?�￰#�����!��6�w�(� �>�0=���P�H��u��u��u����Ï�5߫�N�	'�� � ��I� �  ��
�t�:�È��È�=���Q��� <��� �� � �e���?���ҁI�p�~�e������@!�p@��a�@��@��@���C��C� �T� ��B��C��d��@�7�����3�����K�L�����I�@�m��D�՚��� ����(
%���:T�<�=�x?�ffd�K/]/�C ���/�+R�8��<�/�*>��=�� I���&��6)����<��_>���A!E��<2�!<"7��<L��<`N�<D��<��,0-�j?y/�����"�I�?fff?m?y&�0q�@T싹1�?�`?Uȩ?X��1T��1 ������?��O�7�� |/QO<OuO`O�O�O�O��O�O�O�O_T��5FZ_S__w_�?�_�Ij_�_fXHmN �H[���G� F���_oo
oCo .ogoRo�ovo�o�o�o �o�et}�o`��_T �_{�o����t? ���/��S�>�w��b�U��Uɲ�C@q�֏m����������D�/�T�ç��¬����BH� �� �T��� ������@�I�Y�@n��@��@: �@l��?٧]��� ��%��n�߱���=�=D��������@�o�A�&{C/� �@�U���+J�8��
H��>���=3H���_E� F�6��G��E�A5�F�ĮE���m����fG���E��+E���EX����>�\�G�ZE��M�F�lD�
�п���
���.�� R�=�v�a�������п ����߿��<�'�L� r�]ϖρϺϥ����� �����8�#�\�G߀� kߤߏߴ��������� "��F�1�j�U�g�� ������������� B�-�f�Q���u����� ��������,P ;t_����� ��:%7pz+�(-�4�t�-1���]3����+q4 �{x��+q�0+#����jb/+/1?E�䴛|�0G+ E)�/s/�/�/�/�,.u%Pe2P�.q(?�{4?^?I?�?m9F � �?�?�?�?�?�?�?+r$OOLO7OpO[O�O@;?�O�O�O�Le�O��O1__A_g_U_1)m__�_�_�_�_�_�j  2 H��6+vH�@",c\�b+vB����~�Bȓ�
��A+p@��so+pw�@�o�o�o�o�o-z#o@5o,>P`|k���Tk�k��A8otck�
 `� �����&�8�J��\�n�������#�rr����H-��$�MR_CABLE� 2��( �V`2T0aa@�k�?w��ab���{�?`B?`C �k�O�M�`B���M��.�t D�hr�k����b`�N`By�S`�O
�v7��A��t D�CUkA%W�i�Z`�b`�CW`9-���΋��(ArrD�Q�Z`���*!��S`r �C�/�7 7������|�cD������Z�+u� M�_�į��ͯ����� ݯ�T�O�%�q�I�[� ���ɿ7��!��� (�:�(�i�{ύ�(w*��** ݃�OM �����HV",%�% 234567O8901���� ��P��  � ba �!
כ�n�ot sent ��?�W�%T�ESTFECSA�LGRPg0*badȯԈqF�
��0�0k~h�����(�9UD1:\m�aintenances.xml��_�  �z�DEFAULT�l~݂GRP 2��ʏ  p�tg% � �%1st �mechanic�al checkl�!�������U� �j7�I�[��m��"��cont?roller��������T(���!3E��M��m""8� ���U������P
AC��3�W��@�������C���ge��. battery�G/�U	tI/[/m//�/���Supply greasQ�/�����#<���!�/�U8/??1?C?U?��=�cabl�/�/�?,(
�/�?�?�?O�O�����?�?���?�O�O�O�O�O��$ �O_Ը׿4_ �OY_ k_}_�_�_�O�__&_ 8_�_o1oCoUogo�_ �o�_�_�_�o�o�o	 jo�oQ�o@�o� ����0��f ;��_�q�������� ˏ�,��P�%�7�I� [�m��������ǟ� ����!�3���W��� ����ܟ��ïկ��� H��l�~�S���w��� ��������2�D�� h�=�O�a�sυ�Կ�� ��
������'�9� Kߚ�o߾����Ϸ��� ������N߶�5��$� ��}��������� ��J��n�C�U�g�y� ����������4�	 -?Q��u���� ������f ;��q���� ��,/Pb7/� [/m//�/�/��// (/�/L/!?3?E?W?i? �/�?�/�/ ?�?�?�? OO/O~?SO�?�?�? �O�O�O�O�O2O�O_ hO_�Oa_s_�_�_�_ �O�_�_._oR_'o9o Ko]ooo�_�o�_�_�o o�o�o#5�l�b	 TCp���o ������!�3� E�W�i�{�������Ï Տ�����/�A�S� e�w���������џ������+�=�  }��a?�  @�q �x������v�d�ɯۯ�x*�** �a�f��?� A�S�e�'������������o�c$�¿� "�4���X�j�|�ƿؿ �P�������D��0� B�Tߞϰ�ߜ߮��� 
ߔ�����d�v߈� &�t���Z�������*�<�j�$MR_HIST 2��e};�� 
 \�b�$ 2345678901K�S���J�9�o����s��� �o(����^p �9K����  �$6�Z~� G�k���/� 2/D/�h//�/�/U/��/ �SKCFMA�P  �e�>����p�p��/�%ONREL � �t;��!� �"E�XCFENB%7
8�#�%>1FNCE?74�JOGOVLIM�%7d;�0�"KEY�%7�5�5_PA�N$8�2�2�"RUN�<�5�3SFSP�DTYPe805�#S�IGN%?74T1M�OT�?41�"_C�E_GRP 1��e�#C�[p���O �s|O�O&D�O�O�O_ _�O>_�ON_t_+_�_ O_�_�_�_�_o�_(o �_Lo^oEo�o9o�o�o �o�o�o�o�o6�k��!QZ_EDIT�"D�'CTCOM_�CFG 1��-�H5��� 
vq_/ARC_B2%Ep9�T_MN_MOD�E"F�P9UAP�_CPL�T4NO�CHECK ?^�+ �/ S� e�w���������я� ����+�=�O�a�;�NO_WAIT_�L!GkwV@NT~qѩ�+�ez#��_E�RR`A2��)�!� ��
��.���1S�e�Ԏ��pOᓫ�| �^+qB��B�QW�ڲ��B���jY/���x)<�0�� ?�k�Яk�0���ڒPARAM⒬.�+�O�+R�p'x�!p��� = �� ��������ۿ�ɿ���#�5��Y�k�G�'w��ϯ�B���BOD�RDSP�s$FP8O�FFSET_CAqRap$�	�DIS���S_A�pARK�"GlyOPEN_FILE5�$A�qlv�p�OPTION_I�O�?�1��M_PR�G %�*%$*�����i�WOU��fGP���	�z$��   0� ��z$#���#�	 �hx(#�z&������RG_DSBL  3��!̚����RIENTTO$0�z!C�0�!A ���UT_SIM_ED���"P���V��?LCT ���hr��q�z%d��_P�EX �8�+�RAT� � dP5+��UOP ���|��Б�����z ���z z 2�1���$��2_C�L�X�L�x�� %���+=Oas ������� '9K]o�z'2�����
/ /./@/R/ã�|/�/ �/�/�/�/�/�/??0?B?�il&k/|>��|?�?ϒP�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�?�?_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo�O �OTofoxo�o�o�o�o �o�o�o,>P0b��Coe����}!�����~�����}�}��W�B�{�.� 9�p���������ҏ؏ ���n���<�K�I�p��	`��~�������:�o����ҟ���>o�A�  �e�U'��.����a�k�e?b �������e���q� �������˯��������Os�1� �_� � ��l�@ �]��G�� @D�  Z�?��`�F�?��b���D�  Ez|�9���  ;�	lr�	� �@� 0g��h��� �V�� �� �&�ѱ��H�0#H��G��9G�ģG?�	{Gkf���`S��,���C����\���D	� DO@ D��	�������  �5��>t�[�ù�b�t��� B��Bp�{�!����CO�^���8��� &�`��������6�V��:�(:��:���]�T���p��	'�� � ��I�� �  �<��=��Ͳ���~^��� <���� � ?� �*�^��u�^��5���N���\�&���t�?���C&��C����B[����J���i0]��@�������~�����������
�@��2�v� ��_�\�G���k�����`����������:!����x?�ff0%�"�� [�W�i��8���
>����n���IкX�����������$�>��
�<2�!�<"7�<L���<`N<D��<��,�/>`����
�?ff�f?2�?&l�@�T�~?�`�?Uȩ?X� ��9��gs���b�� `��P��A//:/ %/^/I/�/m/�/�/�/ �/�/�/?�/6?����/?�?+8HmN �H[���G� F���?�?�?�?O �?,OOPO;OtO_OqO �O�E9��M�O%�S?_ w?@_�Od_v_�_�_9 �_�_[_�_�_oo<o�'o���fb�wkC�6o�o2o�o�m?����o�o	�o��çRs��sm��H����Z�d��`�a�q�@I܊�@n��@��@:� @l��?٧�]j ��%��n�߱����=�=D�����p��@��oA�&{C/�� @�U� ��+J8��
H���>��=3H���_
� F��6�G��E��A5F�ĮE���2�D���f�G��E��+�E��EX��Z�D�>\�G�Z�E�M�F�lD�
[���iϏ ���ޏ��;�&�_� J�\���������ݟȟ ���7�"�[�F�� j�����ǯ��į��� !��E�0�i�T�y��� ��ÿ���ҿ���/� �,�e�Pω�tϭϘ� �ϼ������+��O� :�s�^ߗ߂ߔ��߸� ����� �9�$�I�o� Z��~��������������5��r(�q43�9����j�"��3�ϩZ�l��q4� �{�����q�0�+#������jb�����1E�䴛|[
	J8n\(���EP*P��A�O�@��#G2 �MT�x����r$��/� 5/ /Y/ �O�/z/�/�,e�/�/�/�/?,??�A)2?D?z?h?�?�?�?�:  2 oH�6�vH��3\��vBoacao`SB�XpWpA�p@so 8OJO\OnO�O�O�M�CP/�O�O�O__%\U�vN$�p�p�A4T�3�u
  %__�_�_�_�_�_�_ �_o!o3oEoWoio�z�7R����H-���$PARAM_MENU ?
��  �MNUTOOLNUM[1�w��`F�`�`�iAWEPCR�`�.$INCH_R�ATE�`SHE�LL_CFG.$JOB_BASp� WVWPR�.$CENTER�_RIr�`$tAZ�IMUTH OP�TB�a$tELE�VATION T�C�a$tDWqT�YPE SNqA�RCLINK_A�T(pSTATUS��c�y__VALU�q�`LEP�a.$WP_�`�b��| �����$�6�_��Z�l�~����aSSR�EL_ID  �����USE_PROG %�j�%�����CCRT�Ƅ��c�_HOSoT !�j! �]��T� '�y�@�R��{����_TIM�EOU$��g  ~�`GDEBUGƀ��k��GINP_F�LMSKޟ�TRl��PG�p  ���OL�CH��yr
�k�@����ү�� ����C�>�P�b��� ������ӿο��� �(�:�c�^�pςϫ� �ϸ������� ��;��6�H�Z߃��WOR�D ?	�k
 �	RS;�ZPyN�q[MAIpf��SUNq��TE��>ZSTYL5r�ЇCOLX�
��LV�  �U�0��d�TRACEC�TL 1�
n�a � Q ���I�DT Q�
���d�D � ޴��j�������� 7P��UP��p���MP��IP������������	��
��U���
����������0�B�T�������Ȁ Z�l���� �����������@@�@@@@�@@@@ 0	&8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO�bOtO�O�O�O�MI�L1Epȁ]P�`�=�~I�_UP ���[PY��q ���NQY��}d�bG_zj؟�zj�&�_D�EFSPD ���k2Ђ  ���`INPTRL �����a8dU�QPE_CONFIP�X��̈́}aw .$�LIDS��� ~	gLLB 1�X��m��dTB�  B4Vc}fn�Oblj�io�eW_ << ρ?��k�o�o �o�o �o6N lRd�����ZZo��=�4�a��f�Q�C�����ď
eGRoP 1�;l�,��@�  �[��_aA?x�D P��DV�C2���k��E�d-�=��Qw }���o&aY�#´��r�[�B�����������П����_a>'oY>a����K�]�G� =N�=R�b���^��� ѯ�����z��=� �xM�s�^�  Dz����_`
��ɿx�ٿ�� �#��G�2�k�VϏ� zό��ϰ������j��)Q
V7.1�0beta1_d�N B(�A�?\)A�G���F��>��^����F�A���n�f�fF�A�p��AaG��q�q@�����V� ߳�������_cAp@�
�U` �#�5�G�BҢQ�� ���z��v�����`F�B�ga���Ru0��e:��@+�a��QG�@������ B{PB���z�BH�����0�� ��g��;Q*)���x��xR� N�0n��P� �R{�w���W��qdKNOW_M�  �e+VdSV� ����U��I[m��@|��_b5�
cMރ���`�V�	BU���3/�~CT���?��@{Q{�{Pr%n/�,��paMRރ��T��כּ
��/�+̍OADBANFWD��+cSTށ1 1�Y84�Uk�V� l?_VT?f?x?�?�?�? �?�?�?�?;OO,OqO PObO�O�O�O�O�O�O _�O__572@<	!S?_`�<}_Q_߀A3g_y_�_�_574�_�_�_�_575oo1oCo576`oro�o�o57A7�o�o�o�o578�*<57MA 0�6�ds�WOVLD  \{,/ȏ72�PARNUM  �C;��63SCH�y �u
B��P�.3b�UPD��um�|���U_CMP_���p��/',5ĄE�R_CHK҅���,1"�Ϗ�RS8� #?�_MO ?C��_0��U_RES_G?0�\{
��]�� ���֟���+��0� a�T���x���������fP����Я���P� ����`,�K�P��� _`k��������`��ɿ ο��p��υ�Xp�(�G�Lυ�V 1��F�P	!@[l��F�THR_INRп �q�,5d��MA�SS�� Z��MN�����MON_QU?EUE �\u,6TS���TNɀU�qN
�3�J�ENDO�m�i�EXEx�iՎ��BEw�Y�J�OPT�IOV�v�M�PROGRAM %-��%LІ�1�K�TA�SK_I�t��OCFG �-��!�^T�DATA��]�~��2%���� �������/�A�S�e��w�"�����������IWNFO�ǡ�<� ��*<N`r�� �����& 8J\n������ȡ� ��S�I�K�_W��]��ECNB�p�[Q&2/�(GW�2�� �X,		�=����j/�%�!$�N0��)�)���_E?DIT �]��/|�/P�WERFL�����23RGADJ {��*A�  55�?��A5��6M����\u�?�O  Bz3W��<�!���%n�?8�/W3f�2�c7�	HDХl����p1?� A�x��t$F*z%@/'B **:0B ��#O5CQM\ujBeE#��AoI���?�� �O]M�MmOO�O�O�O /_�O�O__!_�_E_ W_�_{_�_o�_�_�_ �_�_soo/o]oSoeo �o�o�o�o�o�oK�o 5+=�as� ��#������ ��9�K�y�o������� ���ۏ�g��#�Q� G�Y�ӟ}�������ş ?����)��1���U� g����������ӯ� ��	���-�?�m�c�u��￙���ٿϿῦ�	 p�zϵ0hϡό�I�πC���ϋ��&�S7P?REF �c:�0��0
5IORI�TY���&�1MP�DSP��:���U�T?�C6ODUC-T<��*)��6;OG�_TG0A���*��HIBIT_�DO	8�TOEN�T 1��+ (�!AF_INE���^�7!tc�pi��!ud����!icmX��>��XY\3��,;��1)� =A�/��0��X�;�G� ��k����������� ��&8\C��	*��\3�c9��?����3>5H�7�B=G/GL�9�4��8��>A�2,  �Y������5
�6)Z)�
//�./�3�ENHA?NCE ճ�2A�d(�/u%��B���J�\�11PO�RT_NUM���0x�1_CARTREP���S2�SKSTA��+�S�LGS[������3�0Unothing�/s?�?�?��<Y?�?�?�?��61T?EMP ����?�8��0_a_seiban��bO��rO �O�O�O�O�O�O_�O (__%_^_I_�_m_�_ �_�_�_�_ o�_$oo Ho3oloWo�o{o�o�o �o�o�o�o2B hS�w���� ���.��R�=�v� a�������Џ���ߏ���<�'�`�O61VOERSI������� disab�le�"KSAVE� ���	26�70H755J�]���!~/�����/�C 	S���:�I�|��e��¯ԯ���J�A��.�9����_��W 1���|��T�ņ����;�UR�GEM B �$���WAFİ ��h"��WW��崖��*WRUP_�DELAY ��>صR_HOT �%_Ƹ�}/e���R_NORMALD����Tϩ�x�SEMI��Ϯ���9�QSKI%Pd�ܺ'u�x[�2� W�V�h�z�=�Gš߯� �������߹���'� M�_�q�7������ �������7�I�[� !��m����������� ����!3EU{�i���G��$R�BTIF�
<RC_VTMOU75��� DCRd�޾� �I�A��3�B�/lB�3�@��M@�7�*�=�������~��� {���T ���j�E��=ߍ�� <2��!<"7�<L���<`N<D��<��,�V���- /)/;/ M/_/q/�/�/�/�/�/��/�/��RDIO_TYPE  k����/EDPROT_CFG ���2��BHͳE�E9
�2�W; ��B�j0�?�:��? ��?�?OM�?KO�� rO�ߓO��O�O�O�O �O_�O5_CWaOf_� -_�_}_�_�_�_�_�_ �_�_1oS_Xow_yoo �o�o�o�o�o�o�o =oBaou�� ������9>� ]��_��������� ݏˏ�#�(�:���[� ���m�������ٟǟ ���$�C��W�E�{� i�����ï��ӯ	�/�� ��G7INT 2��Gɔ1�AG;�� ^�p��2���
Hf�0 ��Ȼ��ٯ �����B�0�f�L�v� �ϊ��Ϯ�������� �>�,�b�t�Zߘ߆� �ߪ���������:� (�^�p�V������������ �6��E�FPOS1 1�~9  x� )c3��������*�w� ����$H��l �+��a�� �2D��+�w �K�o���./ �R/�v//�/�/G/ Y/�/�/�/?�/<?�/ `?�/]?�?1?�?U?�? y?OO�?�?�?\OGO �OO�O?O�OcO�O�O �O"_�OF_�Oj_|__ )_c_�_�_�_�_o�_ 0o�_-ofoo�o%o�o Io�o�oo�o�o, P�ot�3�� i����:�L�� �3������S�܏w�  �����6�яZ���~� �����O�a������  ���D�ߟh��e��� 9�¯]�毁�
���� ɯ�d�O���#���G� пk�Ϳϡ�*�ſN� �rτ��1�k��Ϸ� �ϋ�߯�8���5�n�<�Z�2 1�f�� "�\��������"�� F���C�|���;��� _��������B�-� f����%���I����� ���,��P���� I���i�� �L�p� /�Sew�/� 6/�Z/�~//{/�/ O/�/s/�/�/ ?�/�/ �/?z?e?�?9?�?]? �?�?�?O�?@O�?dO �?�O#O5OGO�O�O�O _�O*_�ON_�OK_�_ _�_C_�_g_�_�_�_ �_�_Jo5ono	o�o-o �oQo�o�o�o�o4 �oX�oQ�� �q�����T� �x����7���[�m� �����>�ُb��� ��!�����W���{�� ��(�ß՟�!���m� ��A�ʯe���$� ��H��l����v߈�3 1��=�O��� ��+�1�O��s�� pϩ�D���h��ό�� �������o�Zߓ�.� ��R���v�����5� ��Y���}��*�<�v� ����������C��� @�y����8���\��� ��������?*c�� �"�F��| �)�M��F ���f��/� /I/�m//�/,/�/ P/b/t/�/?�/3?�/ W?�/{??x?�?L?�? p?�?�?O�?�?�?O wObO�O6O�OZO�O~O �O_�O=_�Oa_�O�_  _2_D_~_�_�_o�_ 'o�_Ko�_Ho�oo�o @o�odo�o�o�o�o�o G2k�*�N �����1��U� ���N�����ӏn� ��������Q��u�����4�������4 1���j�|���4�� X�^�|����;���֯ q��������B�ݯ� �;�������[��� ϣ��>�ٿb����� !Ϫ�E�W�iϣ���� (���L���p��mߦ� A���e��߉��߿� ���l�W��+��O� ��s������2���V� ��z��'�9�s����� ������@��=v �5�Y�}� ��<'`�� �C��y/�&/ �J/��	/C/�/�/ �/c/�/�/?�/?F? �/j??�?)?�?M?_? q?�?O�?0O�?TO�? xOOuO�OIO�OmO�O �O_�O�O�O_t___ �_3_�_W_�_{_�_o �_:o�_^o�_�oo/o Ao{o�o�o �o$�o H�oE~�=��a�П�5 1� ퟗ��a�L���� ��D�͏h�ʏ���'� K��o�
��.�h� ɟ��퟈����5�П 2�k����*���N�ׯ r�����Я1��U�� y����8���ӿn��� ��϶�?�ڿ���8� �τϽ�X���|�ߠ� �;���_��σ�ߧ� B�T�fߠ����%��� I���m��j��>��� b����������� i�T���(���L���p� ����/��S��w $6p���� �=�:s� 2�V�z��� 9/$/]/��//�/@/ �/�/v/�/�/#?�/G? �/�/?@?�?�?�?`? �?�?O�?
OCO�?gO O�O&O�OJO\OnO�O 	_�O-_�OQ_�Ou__ r_�_F_�_j_�_�_o<��6 1���_ �_o�oyo�o�_�oqo �o�o�o0�oT�ox �7I[��� ��>��b��_��� 3���W���{������ Ï��^�I������A� ʟe�ǟ ���$���H� �l���+�e�Ư�� ꯅ����2�ͯ/�h� ���'���K�Կo��� ��Ϳ.��R��v�� ��5ϗ���k��Ϗ�� ��<�������5ߖ߁� ��U���y�����8� ��\��߀���?�Q� c������"���F��� j��g���;���_��� ��������fQ �%�I�m� �,�P�t! 3m����/� :/�7/p//�///�/ S/�/w/�/�/�/6?!? Z?�/~??�?=?�?�? s?�?�? O�?DO*o<d7 1�Go�?O=O �O�O�O�?_�O'_�O $_]_�O�__�_@_�_ d_v_�_�_#ooGo�_ koo�o*o�o�o`o�o �o�o1�o�o�o* �v�J�n�� �-��Q��u���� 4�F�X����ޏ��� ;�֏_���\���0��� T�ݟx���������� [�F�����>�ǯb� į����!���E��i� ��(�b�ÿ��翂� Ϧ�/�ʿ,�e� ω� $ϭ�H���l�~ϐ��� +��O���s�ߗ�2� ����h��ߌ���9� ������2��~��R� ��v������5���Y� ��}����<�N�`��� ������C��g d�8�\��	 ���cN�" �F�j�/�)/��M/�q/WOiD8 1�tO/0/j/�/�/ ?/0?�/T?�/Q?�? %?�?I?�?m?�?�?�? �?�?PO;OtOO�O3O �OWO�O�O�O_�O:_ �O^_�O__W_�_�_ �_w_ o�_$o�_!oZo �_~oo�o=o�oaoso �o�o D�oh �'��]��
� �.����'���s� ��G�Џk�􏏏�*� ŏN��r����1�C� U����۟���8�ӟ \���Y���-���Q�گ u�����������X�C� |����;�Ŀ_����� ��Ϲ�B�ݿf��� %�_��ϫ����ߣ� ,���)�b��φ�!ߪ� E���i�{ߍ���(�� L���p���/���� e�������6����� ��/���{���O���s� ������2��V��z���/�$MASKW 1�+�����XNO  ����MOTE � �$G_CFG� �N��P?L_RANGJ?��%��OWER ��%��SM�_DRYPRG %�)�%K��TART ��	*UME_PRO���e/�$_EXE�C_ENB  z?�GSPD> � �(�(TDḄ/�*RM�/�(IA_OPTION����!_A�IRPUR� pF*B?�MT_� �T�L�`1g��o=�"C�?  N?�?�?�?�??1�OBOT_ISO�LC�>0~z�ENAME �F*T/�	OB_C�ATEG� ��O�DuCORD_�NUM ?��;1H755  ?�O�OY� �PC_TIMEO�UT� x� S2�32g1��#� LTEAC�H PENDAN0!Pc�pT�=J�H Mainte�nance CoKns?m_?"�_�DNo Use �=�__�_�_oo%o�9RNPO #R��56QCH_LfA �?� 	�a~so!UD1:�ozuoR� VAIL�A�5�1SR + /;1��e�R_INTVAL�6��Yp> yV�_DATA_GR�P 2�� D>pP��� ��y�!��A�/� e�S���w�������� я���+��O�=�_� ��s�����͟���ߟ ���K�9�o�]��� ������ǯ�ۯ��� 5�#�Y�G�i�k�}��� ��׿ſ�����/� U�C�y�gϝϋ��ϯ� �������	�?�-�c� Q߇�uߗ߽߫�����$SAF_DO_PULSK�A? <��CSCANR6��<@SC�� �`!X�!�? �1
@�2��A�Q�U[�? ����������� |��#�5�G�Y�k�H+rc�2��[�"��d����>	X�Hi @�����?���. �p�/_ @3T01�n���YT D������� "4FXj|�������BoLe���V,/>/F$�
*  iU;��o�Tg!EqpduE
�t��Di�@��k�Z  � �+Jk���AS��/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_.a����_�_�_oo)o ;oMo_o�_���o�o�o �o�o�o�o	-2qoo0�"�#�%�-~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�N� �_r���������̯ޯ ���o8�J�\�n� ��������ȿ3auk ���,�>�P�b�t� �ϘϪϼ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{��������(������ /�A�S�e�w������� ��������+=���
�T�������"z�	12345678�"�h!B!�Q��������f� �'9K]o ��	������ //(/:/L/^/p/�/ �/�/�/�/�-��/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO�/ �/TOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_3O�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�_�o  $6HZl~� ������� � �oD�V�h�z������� ԏ���
��.�@� R�d�v�5�������П �����*�<�N�`� r���������̯��� ��&�8�J�\�n��� ������ȿڿ����D"����D�V���{ύϟϻ
Cz � Bp��   ����2�� _} 6��
�ǿ�  	���2@<�#�5�G�Y�i���j��߯��������� 	��-�?�Q�c�u�� ������������� )�;�M�_�q������� ��������%7@I[m��� j��k����<� ���  �������
�
�t�  ��
"��`��$SCR_GR�P 1�!*P�!30� � }��� ���	 m�u�k�����ǒ�����ٰ���C� ���݌*'���L�R Mate 2�00iD 567�890�LRM�c# 	LR2D� j ��
123�4i%�x�m�� �&_u��d�d��ӻ����)	��"?%?7?I?[?k<��H�u�$yd�?��?�?�?�#����?(O�?LO��>K� h��,W���eEB���Ɛ�O�B�D�A���O c @���E�@��@F�O ? �E�BH���_�J�F@ F�`8R@_7Od_O_�_ s_�_�_�_�_�_o� �A�AR1oo.o@oRdB�`o�_�o�o�o�o �o�o�o$H3l W�~ߥz#��w�����������A@� >��,��@h�@U����k��' �,�;ϫ���A�@�vH΅�?�5ۀ���"��� ��*��z��M�Y�k�:�h���
 ����ß��ҟ����Y/k#DECL�VL  ������"܂A��*S�YSTEM*��V�9.10214 �s�8/21/20�20 A � �`�o�SERVE�NT_T   �$ $S_NA�ME !��P�ORT����RO�TO�� ��_SP-D��J�B�̠�TRQ   �
ɣAXISҡ�קϠ 2 �ɣD�ETAIL_ � l $DA�TETI����ER�R_COD(�IM�P_VEL�� �	:�TOQB�AN�GLESB�DIS蜠N���G��%$L�IN(� ȤREC�ҡ ,�����F�MRA�� 2w d��IDX��܋�ߠ h�$�OVER_LIM�I��栄0ɣOCC�URҡ  �-�COUNTER������SFZN�_CFGҡ 4� $ENABL�(�ST"���FLA�G��DEBUF�R�[�J��Jҡ �� 
$MIN_OwVRD��$I���W�{�s���FACE��|�SAF��MI�XED�̄�d�{�R{OB��$NE��{PPôHELL ��	 5$J���BAS(�RSR�_.�  $N�UM_�B� R�1w��29�39�U49�59�69�79�98w�	�ROO��~�{CO��ONLY�p�$USE_AB����ACKEN�BA���IN۰T_�CHK��OP_S�EL_9���_PUl���M_%�OU��PNSֽ���x�9����M3�TPFWD�_KAR@���.�R�E��$OPTI{ONX�$QUE �꿠D;�Y��$CSTOPI_AL�ӆ��EX���ь�(�X�T��M1��2��M�A��STY��SO���NB��DI��T�RIFÄ�@�INIr��Mà��NRQ���END��$K�EYSWITCH�'�<����HE=�B�EATMo�PEROM_LE?�G�E<�Jn�U;�F��<�S��DO_HOM��O����EFP����Gæ�STL��C��O�M)���OV_MS��ѻ�ET_IOC#MN�Ӕ���]����HK��
 D �-Ǳ�SU'���MP���.�PO��$F�ORC&�WARNvOM� �@?$FUNC� 7ÙU���AR���2j�3�4~ �*�OL�Lo��!�OUNLO�%���ED%��p�SN�PX_AS#� �0$�ADDV�X��$SIZ(�$V�ARw�MULTI�P���� Ao? � $�� ���	&�� ��'�C<;�kFRIF��۰aSl�~	��[NF��ODBUS_AD`�&ү���CM1��DIA]$DUOMMY1���3��4��SО� g� X�TE���8�SGL#!T}A��  &8��<#'�� 5 $ STMyT��U#PSEG���U!BW��%$SHO�W]%��BANi T�POF��9�0����ȠVC��Gvh� 1 $PC�ܰ� �$FBkP�(SP��A���%��VD� g�� � �A0��0�b� $1� +7� +7� +7� �+75)96)97)98*)99)9A)9B)9}  +7�+7r +7F)8�  �859��8O9	 �8i9U1v91�91�91�9U1�91�91�91�9�1�91�9���G592�B92O92\92i92�v92�92�92�92��92�92�92�92��92�93(93593�B93O93\93i93�v93�93�93�93��93�93�93�93��93�94(94594�B94O94\94i94�v94�94�94�94��94�94�94�94��94�95(95595�B95O95\95i95�v95�95�95�95��95�95�95�95��95�96(96596�B96O96\96i96�v96�96�96�96��96�96�96�96��96�97(97597�B97O97\97i97�v97c�7�97�97��97�97�97�97��97�42 � Pzk�UТ ٠Ĩ�.�
1��� x $TORu�V�  D�M��RΠ,��ߔQ_��R��P�(�G B�S��C=���'�_U� 2��Y�SLu��� � �3ǚ
J�$0x��^��"VALU3����A�����FO�ID�_L���HI��I~]$FILE_����$��7M�S=Aϱ hҐ�?E_BLCKo�#�|>!,�D_CPU<��<�
>����ǰY�# �R  � PW���В��LAc!Sα�������RUN_FLG ŵ��ɱ��?�̵걡�걬�Hิ���b�T2A�_LIo�  �G_O���I�P_EDI���0T2��,��4��	��7�]�@��TBC24 �� ��̰� ��,�FqT�����TDC̰A��C���M�����&��TH�S������R��� . ERVAE�������������� X ;-$:�LEN��G���:в�RAk��N��W_�i�1:�פ2&��MO4��S���I��#�㡩�Ք:о��DE�աLACE����CC�#��_�MA� ������T#CV�/���T!�0� O�E�2���!s����!�J��A�%M�䟠JH�0������Fс2���0����� JK��VK�!���������J�!���JJv�JJ�AAL��@1��1�+�
!/�5��b�N1V�b�!��!��L��_Q!������C�F� `ҐGRCOU��?!��!N���CS��REQUI9R�EBUj6�n��$T��2���7������ �� \�w f�APPR��C�L!�
$=�N0CLOr�@	S��U	�չ
��> �n�M����a���_MG�� C0��0	��BRK�	NOLyD�� RTMO+�H�
��J+��P3� ��������O���X�J��6 7 1!H�|6ц�� ���a��!���PATH����f؟� ��%�� SCA�j��1�IN9�U�C�Д��C0UM(Y������	!á��$*�$*:$ PA�YLOA�J2L���R_AN��e#L���o)k!_){!�R_?F2LSHR	Ԩ!LOp$��'#�'#ACRL_y��� ��W$�H��!�$yH�2FLEX3���J�� P��ϧ�� ߞ�#�B}J9�  :F� X��Щ7�4[����d�v߈�F1�1E"G��@�߻�������RBE�� ��1�C�U�g�y�� )XFT�����6@XX����1��T�W'QX �0Q��D}H���U�H ����0�4�=�+�O�`X�j�|���"�BJ��! �����������Ƭ�AT;F���ELP�@�s��J�� ��;JE� CTR�6A�TNƑ	v��HAN/D_VB!�31��nt" $�PF2�����SW��2�~#� $$M�  �	���x��|�@�u�vAƠ\ �š���A����
A�A����U��
D�D��P�G����ST�����	��N�DY ˰. ��t�} ;П' �1�'�!^'��}T�0�P�P(1:CLU�^gyJ��$ �p�4� cA��b���ASYM�#�����#���!�_ ��(�$����x/-/?/Q/c#Jj,|*p�����)HD_VIds�٨b�V_UN K�ؠ�� c�!J��� E���,��%(�L��-����)�/?���S0$4,3l��HRt�i��%zrͱF0@�DI� ��O���ΰ�c�& 0`�I�A �#�<@'�'�?@|����Aϰ ' �� �qME�A�t`B�)�T�PT@��`�j����E0�a�oȊ�~�T����� $DUMMY}1:$PS_9@�RF�0  ���n� FLA��YP�S���r�$GLB_T�p���j�N1�0x@:qF�( X ��t�ST�A��SBR��M21_V��T�$SV_ER� O���@�X�CL�@�A��@O�ɰGL�E�W��) 4��t�+$Y!bZ!bW������!�sAC�"����U.��* �PN�Ѕ��$GIJp}$>�� )x�ӼЎ��+ L����S�}�$FS�E��NEA�R�@N@CF-�@T�ANC@B��JOG��0 ,�0$�JOINT�Q�P� ��MSET��-�  ��E�A�`S��bjp���`��.�k BpU�A?���LOCK_FO� ��q�BGLV=sG�L��TEST_X9M3 ��EMPi���q�����$U�0����P2*���!�+���p��!�)B�CE�����B� $KAR��AM�TPDRA8��_�V�VEC�0p��Z�IU!�,&�HE���TOOLC��VvDREw�IS3�5r��6C6@ACH|����-��O�rô�3�0a��SI# � @$RAIL_�BOXE�Qe�R�OBO��?�e�HOWWAR1����ROLM��7�a���H�a��*@vO_�F�`!e�HTML5��������Rw/b�mRz�O�2�0b��0k�o ��O�U~�1 d���)�)�r�a��$PIP��N�P������H@�!� �0CORDEaD���� *�XT� ���)ɰ�`O)� �2 D ��OB E�s��P?����?�S�qSYS?ADqRqɰj�TCH�p� 3 ,�PENTҲO1A��_�����a'��PVWVA~E�4 � e�����PREV_R�TR�$EDIT��VSHWR�aP,� �B��٠DT��1'$ a$HECADd���A t���KE�Ѩ�CPSP]DX&JMP\L��R�TR�@�5�GD1�I��SrC�^pNE��qTwTISCKC�MM1�q��#HN"�6 @pI�!�e`!_GP�&���P0STY���L�O��ӂ"�"�07 �t 
�G�%$����=,�S`!�$��PY������P��&SQUY��5��ءTERCn�!a��=S�d8 ��8�@�g�P�g%Q���`Oo��b�D@IZ��������PR%��B�!� sPU�aE_DO2�֫XSz�K�AXiI<@[&�UR�`��Cr � j�q�`_,��|ET}BP��X ҕ��d Ӗ<0A߁Ց��9��)����{SRqt9l�0 �y�R�z�E�v
Y�r�E �w�C��C�>U3�>U C�>US�PUj]��PU�\$��nYC�_|]C�]L�p^�p����qSSC��� : he�DS�� `��SP�jeA	TA��rA� �"�¿ADDRES��B��SHIF�c�_W2CHpfIЮ�a�TU�I�q �;b�CUSTOT�D��V��I�<�P��~aC��
��
�rqV�-AG�= \*Ђ��;0|�1�0IrC���2�Bz�^�Iq�TXSCREEA�>ٰW1TINA�{��Мt����� Q_~b��? T �![�B|Z�7��vJAp{JB�t�RRO��G�{R �qbD�UE��$@ ������S�|�|RSM� @GU`.�0�S�ͰS_�Ӏs��c�v����~ACx��O��t 2?��UE��A�kҶ�@WGMT_�L9�YA�G�Ol����BB�L_��W��G�B ��;0�O���L�E�b*� �b)�RI;GH3�BRDmԤaOCKGR��[�T/|Z�W�WIDTH�� aB������2�I&j EY~`F�C�z �6 2��	ABAC�K1��Εq�M�F�O�LAB(Q?�(M�I����$UAR�S৐S�H	�� D 8��G�_@!�b1�T�R�����C������0�O�aG�E�� x�T�U?��R��BLUM�aF�`�ERV�1�IH�N�E��FK��@GE`��@5I LPѥ�BE�0/a)�?a��POa������5��6��7��8ޢ�2b�@1�]t������S�0�E��USR��G <*�S�U���c��sFO�`��PRI�A�m��m�аTRIP���m�UNDO
�H��`0�BE)�AE��{@u0 qI,���AG H0aT[ a�a'�OSr��<�R�@�Û�ӁJ��ߤӫ�c��$�p�U١ӁKl�~ό�٢�%N�OFF����L(�%��O��"�Je���Z�Ke�GUvP��m��a)׻�SUB8�"t�̀SRTe��DaM�"F�g �3OR��No�RAU�@p�T���U�_��$N |��@�OWN���$SRC���^0Dx�����BMPFI4a}@ESPA�2�p ����.!��������
 nӁO `��WO$Pr��1�0COP��$r@�_�м�i�,�p�WA�C�� M�#�L��� �5�a� P�rSHAD�OW^@���_UN�SCA~�㓔��D�GD��WEGAC<c�w�VC P)�>ӁQ� ��@6l3$�ER�p,�Ȁ1����C� ,�DRkIV�6�A_V� �O�� 6 D|�MY_UBY{�4�B6c�l5��0�p.!��1���P_��4��L#KB�M&�$� DEYƧEX �'�t�MUbv X&�h�USz!h@˰_R�q�2���`���1G�PPACIN�!i0RG��Xn���n��n��i�REF��ac�,��n��R �`[�Gt�P�r� ���RS��S ��x����O�	h�:A�RE+SWf _A$g.� @O���aQA�`'�BEl�U.0dH�-��`�HK32Tu�?�0�A$�ppEA� zL�3�'����MRCVӁU� �ʠO?0M3�Cs	��ð�REF��������C � ���!�!�1%�f_��|g(�xPSi����1{1��ЄV �2�����04�����0OU�'�<�&4� Q�a�2��$�p_p@���S}ca�!D��`UL6�pT(�COG�H�3U 0NT#�P4�1�O5`�[6��[30L���5��5`��7����VIA_L�]`W� ��HD�`Ɛ�$JOg����?$Z_UPL̰ �ZEPW�5�139����_LIM�$EP 1I�4��1�1�q�a���`��0&�6�Xģ 0}c�A@` }cC7ACH��LO!lD@�A �I��|���C@KMI�cFA�ETVP��F�+$HO3����p@COMMJ�O�O =��G�'��d3��͡�$� �VP�p�6R_SIZ��@TZR ;X�1�<W��n�MP`ZFA�I�0Gl�@AD�Yi�MRE�$�REW�GPU� ��s�AS�YNBUFs�VR�TD�U�TEQn�OL��`D_��
eW��PMC�`TU �@QD��UECCU�VE�M� �ERb�GVIR�C�Qe�SN��Q_DELA����簶��AG�YRXYZ��}�W��h!�dd��o`T�IM�a�f�b���EGRAB�B`�Y+�%�ЄY:��ڒLAS��;.PA_GEWEZ>���sbc_uT�#���)�����I�t��fb�BeG/�V��p�PKq X�fXA�'GIOpN쐒)%s�0G�Q:�[$���AS�P}FN�� LEXPv\��ӳ��z�Q��I �S�� E���E���md��b����]��+��DY������F�ORDı���°@��"�^ $.0TIT�ɰ�8�����VSFv��Ӈ_  ��$�[1 U�R��PSM�`����ADJ΀�0;ZD�a D��A�AL�0�PΠ
BPE�RI<@��MSG_Qc$FQdU����eBa�b���0�@��6�@�W�XS�h�Qc��� K�CH)�HOL�� ��X�VR�d7r+�T_�OVR2��ZABC\�e�6��C��
�1c�z�VS@ f � $_�<��|�CTIVz��A�IO���FY�ITl
�mDV	�
m�X@��{Q��àP	S�!�� �S���A� ���ALSTY��A�0l0��_S��MA�c�DCSCH��g Lg�#�w��@ �G�8�@� EPGNA�C��x�A"�_FUN�>�@	 �Z&�촙h���$L������ZMPCF\�i����
�����LN� �.�
���`]�j $�Az���CMCM` Cr�C�\���9P^� '$J��D+Q!� 2�+ǚ07Ś0Ǩ���0�c�UX�a��UXE&���a&�z�<�z�����Ɍ����FTFp<1!���; �Z�k D���4�ٰ��Y@Dp l� 8cR�PU��?$HEIGHv�#?(0ؖ����>�$m � �S��$B0A���L�SH�IFvS��RV@F�����+�C�0�\� -4�D��ְ^s�� UYD���CE��V}!}x��SPHERh� n ,00�F�fX� �r���FA;1���c���u��S�HOT��_��@S�MIP�OWERFL  �c� k�R��W7FDO`� ��G@~� 1 ����ᾌ� L!��_�EIP���c��j/!AFz0E_�$����!FT��S���w�!�x�����f���!R'`MA@����������p��������[!O�PCUA\�
<J�!TPz0p���d��!
P�M��XY��e �?�	�f.�_!RDM�V���gz�!R9�0�	�h�#/!
����@X�i/o/!�RL�PCp/�)�8^/�/!ROS����,�4�/?!
CE� MT�@?�Yk�/S?!	2C{�dq?�lB?�?!2�WASRC��m�?�?!2USB��?�n�?7O!S#TM��QO�o&O�O@���O�tO�M��I
��KL ?%�� �(%SVCPR#G1�OZU2__"P3@_E_P4h_m_"P5�_�_P6�_�_"P7�_�_P8ooP90o5kT�]o Q
_�oQ2_�oQZ_ �oQ�_�oQ�_%Q �_MQ�_uQ"o� QJo�/Qso�/Q�o �/Q�o=�/Q�oe�/Q ��/Q;��/Qcݏ /Q��/Q�-�/Q� U�WQ��O�BG`�O P ���'Q����1�� U�@�y�d�������ӯ �������?�*�Q� u�`����������̿ ���;�&�_�Jσ� nϧϒϹ�������� %��I�4�m��jߣ� ���߲��������!��E�0�i��J_DEV� ���M�C:t��GRP �2��� �@bx� 	� 
 ,��q��﬒����� 9� �2�o�V���z��� ��������#
G .k}��X�� ���1U< y`r����� 	/�-/�"/c//�/ n/�/�/�/�/�/?? �/;?"?_?q?X?�?|? �?�?�?�?F/O%OO IO0OmOTOfO�O�O�O �O�O�O�O!__E_W_ >_{_b_�_�_O�_�_ �_o�_/ooSoeoLo �opo�o�o�o�o�o �o+=$a�_V� N������� 9�K�2�o�V������� ɏ���ԏ�#�zG� Y�@�}�d�������ן ������1��U�<� y���r�����ӯ�<� 	���-�?�&�c�J��� ���������ȿڿ� ��;�"�_�q�Xϕ�� ���ς������%�� I�0�m��fߣߊ��� ��������!���W�.��d �^�	E��y���������	�%��	�.������ G���G�W�e�O���s� ��������� C��� -Q?acu� �����) M;]����� ��/�%//I/� p/�9/�/5/�/�/�/ �/�/!?c/H?�/?{? i?�?�?�?�?�?�?;?  O_?�?SOAOwOeO�O �O�O�OO�O7O�O+_ _O_=_s_a_�_�O�_ �_�_�_�_�_'ooKo 9ooo�_�o�__o�o�o �o�o�o#G�on �o7������ ��aF���y�g� ��������я'�M�� ]���Q�?�u�c����� �����#������'� M�;�q�_���ן���� ���ݯ��#�I�7� m�����ӯ]�ǿ��� ٿ����Eχ�lϫ� 5ϟύ��ϱ������ M�2�D������eߛ� �߿߭���%�
�I��� =�+�M�O�a���� ����!����9�'� I�K�]��������� ������5#E�� �����k���� �1sX�!� �����	/K 0/o�c/Q/�/u/�/ �/�/�/#/?G/�/;? )?_?M?�?q?�?�?�/ �??�?OO7O%O[O IOO�?�O�OoO�OkO �O_�O3_!_W_�O~_ �OG_�_�_�_�_�_o �_/oq_Vo�_o�owo �o�o�o�o�oIo. mo�oaO�s�� �5�E�9�'� ]�K���o����̏� �������5�#�Y�G� }������m�ןş�� ��1��U���|��� E�����ӯ������ -�o�T������u��� ��Ͽ���5��,�� �߿Mσ�qϧϕ��� ���1ϻ�%��5�7� I��mߣ�����	ߓ� ����!��1�3�E�{� �ߢ���k��������� ��-����z���S� ������������[� @�	s��� ���3W�K 9o]��� �/�#//G/5/k/ Y/{/�/��//�/�/ �/??C?1?g?�/�? �?W?y?S?�?�?�?O 	O?O�?fO�?/O�O�O �O�O�O�O�O_YO>_ }O_q___�_�_�_�_ �_�_1_oU_�_Io7o mo[o�oo�o�_o�o -o�o!E3iW ��o��o}�y� ��A�/�e����� U������я��� =��d���-������� ��ߟ͟��W�<�{� �o�]���������ۯ ���˯�ǯ5�k� Y���}�����ڿ��� �����1�g�Uϋ� Ϳ���{�����	��� ��-�cߥϊ���S� �߫���������k� ��b��;����� �����C�(�g���[� ��k�����������  ?���3!WEg �{����� �/SAc�� ��y��/�+/ /O/�v/�/?/a/;/ �/�/�/?�/'?i/N? �/?�?o?�?�?�?�? �?�?A?&Oe?�?YOGO }OkO�O�O�O�OO�O =O�O1__U_C_y_g_ �_�O_�__�_	o�_ -ooQo?ouo�_�o�_ eo�oao�o�o) M�ot�o=��� ����%�gL�� ��m�����Ǐ��׏ ��?�$�c��W�E�{� i�����ß������ ՟���S�A�w�e��� ݟ¯�������� �O�=�s�����ٯc� Ϳ���߿���K� ��rϱ�;ϥϓ��Ϸ� ������S�y�J߉�#� }�kߡߏ��߳���+� �O���C���S�y�g� ��������'��� 	�?�-�O�u�c����� ���������; )Kq�����a� ���7y^ p'I#���� �/Q6/u�i/W/ y/{/�/�/�/�/)/? M/�/A?/?e?S?u?w? �?�??�?%?�?OO =O+OaOOOqO�?�?�O �?�O�O�O__9_'_ ]_�O�_�OM_�_I_�_ �_�_o�_5ow_\o�_ %o�o}o�o�o�o�o�o Oo4so�ogU� y����'�K �?�-�c�Q���u��� �ҏ䏛������;� )�_�M���ŏ���s� ݟ˟���7�%�[� ������K�����ٯǯ ����3�u�Z���#� ��{�����տÿ�;� a�2�q��e�Sω�w� �ϛ������7���+� ��;�a�O߅�sߩ��� ��ߙ����'��7� ]�K���ߨ���q��� ������#��3�Y��� ����I����������� ��a�FX1 y�����9�]g�$SERV�_MAIL  �g]�COUT�PUTR�h @GRV 2��  ` (��-�GSAVE�saTOP10 �2� d  c/+/=/O/a/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O��O�O�O_��YP��DFZN_CF�G ��`$��MQGRP� 2WW� ,�B   A�PgD�;� B�P� � B4#RB{21�HELLPRC	����nW| ok%RSRo o"o[oFoojo�o�o �o�o�o�o�o!E�0i{�~�  �]r����r� h ��r�q�x
�r2h d�|�}8��V�HK 1
�[ �r�|�v���ɏď ֏����0�Y�T��f�x����������\OMM �_��R�FTOV_ENB�R��P�OW_R�EG_UI0�EIMIOFWDL������Ue�WAIT�-�1�oR��mQ�ܚ��TIMQ����įVAQ��e�_�UNIT,����L]CJ�TRYQ���GMON_AL�IAS ?e���he������� úm����
��ǿ@� R�d�vψ�3ϬϾ��� ���ϟ��*�<�N�`� ߄ߖߨߺ�e����� ��&���J�\�n�� ��=����������� "�4�F�X�j������ ����o�����0 ��Tfx��G� ����,>P bs����y �//(/:/�^/p/ �/�/�/Q/�/�/�/ ? ?�/6?H?Z?l??�? �?�?�?�?�?�?O O 2ODO�?hOzO�O�O�O [O�O�O�O
_�O_@_ R_d_v_!_�_�_�_�_ �_�_oo*o<oNo�_ ro�o�o�o�oeo�o�o �o8J\n� +������� "�4�F�X��|����� ��]�Ï�����ɏ B�T�f�x���5����� ҟ������,�>�P� b����������g�� ���(�ӯL�^�p������>��$SMO�N_DEFPRO�G &������ &�*SYSTEM*���߷p��?���RECALL �?}�� ( ��}4xcopy �fr:\*.* �virt:\tm�pback#�=>�169.254.�@�120:450�4 J�S�e�wφ�}5�a"�4�F�P�������}9�s:o�rderfil.dat�̺���a�s����}0�mdb: ��>�K�K����� �� ϬϹ���`�r��π(�:�����������xyzrate 124 �����[��m����!�:�1708��=�O����� }:�,ߥ���Tfx��1��5��L �����5����as�}6��+=� Q���tp?disc 0������\/n/�/��t�pconn 0  ;/5/G/�/�/�/! �EV?h?z?��:? ��?�?�?�A �?dOvO��,O>OQOh�O�O�O
�1 �O �O�OZ_l_~_������ G_�_�_�_?!?�?E? Vohozo�?�?:o�?�o �o�oOO0_AO�od v�O�O,>Q�� �o+o�o�o`�r��� �o2��oM�ޏ��� ���K\�n����$� 6��ڟ����#��� ǟX�j�|�� �_@�964�/L�ݯ�� �&�����S�e�w��� ��7���K�ܿ� �� &�8���Ͽ`�rτϗ� (�:ϸ�P������� �ϼ���_�q߃ߖ���664�/K����� ��/�ٸ���[�m� �/$�6�H������� �"�����S�e�w��� ��7���K����� ���$SNPX_A�SG 2����%� � ��%�M � ?�PARAoM %/� �	;P�r�P��& � OFT_KB_?CFG  �+�OPIN_SI�M  %���( RVN�ORDY_DO � ��:QS�TP_DSB���~SR �%	 � &2 A�B_WELD_1����TOP_ON_ERRG��PTN z% �A	"�RING_PRM��YVCNT_G�P 2��2 x 	zy/�g/�/�/��/VDN RP 1u	� �!%�/ �/?#?5?G?n?k?}? �?�?�?�?�?�?�?O 4O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _o�o�o�o�o�o�o�o �o%LI[m ������� �!�3�E�W�i�{��� ����؏Տ����� /�A�S�e�w������� ��џ�����+�=� d�a�s���������ͯ ߯��*�'�9�K�]� o���������ɿ�� ���#�5�G�Y�k�}� �϶ϳ���������� �1�C�U�|�yߋߝ��������"PRG_�COUNT��"��ENB4/��M�$��1�_UPD �1�T  
 ���{��������� �����/�X�S�e� w��������������� 0+=Oxs� ����� 'PK]o��� �����(/#/5/ G/p/k/}/�/�/�/�/ �/ ?�/??H?C?U? g?�?�?�?�?�?�?�? �? OO-O?OhOcOuO �O�O�O�O�O�O�O_ _@_;_M___�_�_�_ �_�_�_�_�_oo%o���_INFO 1=i�O�q`	 Ho�owo�o�i�?���bf;�>����c�8��o B�B��QW�ڲ�B����jY���ɻo.~ �C��CB���Õ���v2����IBB��L?q�D�B��jA{"Op�SpEC
���Y?SDEBUG	�j���?`dR�zpSP_�PASS	�B?~�{LOG ff]s�  ?`.x�Eo  �N�?aUD1:\�tLn�r_MPC�}i�:�L��i��qj� i��SAV �y�q��q�r;e �SV��TEM_TIM�E 1�wt� 0O�;K�� �;d�ʇMEMBK  i�N��p�N��`�p�X|O��3 @p�;cВ����ǜ�������q {@�/�A�S�e� ��}�������ůׯ� ���!�3�E�W� i�{�������e��ӿ ���	��-�?�Q�c� uχϙϫϽ�������0��)�̅SK%�*���9�i�{ߍ߁�4�?`X,�2����A���p �>b ֒" ��� ��$�T�f�x�<l���  ����Ԁ;c����������߀�+�P�b�t�����?`$ ����������, >Pbt���� ���(:.��T1SVGUNS�PD�u '�u��]2MODE_LIM ,�恐rY�2f��}XA�SK_OPTIO�N�p-��q�_D�I�pENB  ��Ռu�BC2_GRP 2LՌs삘$/Ւ�C�9#QBCCFG +Ƨ� ���/t&` �/�/�/�/�/�/ ? ?D?/?h?S?�?w?�? �?�?�?�?
O�?.OO >OdOOO�OsO�O�O�O �O�O_���L _�OS_ e_�OB_�_�_�_�_�_ q�o/��Po1ooUo Coyogo�o�o�o�o�o �o�o	?-cQ s������� ���)�_�E�0Ps� ������ǏE��ُ�� !��E�W�i�7���{� ����՟ß����/� �S�A�w�e������� ѯ�������=�+� M�O�a�������q�ӿ ���'ϥ�K�9�[� ��oϥϷ��ϗ����� ���5�#�E�G�Yߏ� }߳ߡ���������� 1��U�C�y�g��� ����������ѿ3� E�c�u���������� ����)��M; q_������ �7%[Ik ������� //!/W/E/{/1��/ �/�/�/�/e/?�/? A?/?e?w?�?W?�?�? �?�?�?�?OOOOO =OsOaO�O�O�O�O�O �O�O__9_'_]_K_ m_o_�_�_�_�_�/�_ o#o5oGo�_koYo{o �o�o�o�o�o�o�o 1UCegy� ������	�+� Q�?�u�c��������� ͏Ϗ���;��_S� e�������%�˟��۟ ��%�7�I��m�[� �������ůǯٯ� ��3�!�W�E�{�i��� ����տÿ����� -�/�A�w�eϛ�Q��� ������߅�+��;��a�O߅�o֣��$T�BCSG_GRP� 2o���  �� 
? ?�  ���� �����(��$�^�H�Ђ��Ү���d�@ ���?��	 HBL������?B$  C�����	�����Cz	�Q�A�Д�333?&f�f?����A�����a� ���͘��|���DH����@��q��t� ����D"w�����d/
 ��r����u������:I�c	V3.00~��	lr2dI	*�}�ҔS3 � ���  �/+��J2����fG/$%�CFG !o�e�� ��K*�u"q�x,�,��/ �/�*x��/�/�/?	? B?-?f?Q?�?u?�?�? �?�?�?O�?,OO<O bOMO�OqO�O�O�O�O �O�O�O(__L_7_p_ �_�����_�_�_[_�_ �_�_oo>o)oboMo �o�o�o�owo�o�o �o:�я�_k�o q������� %��5�[�I��m��� ��Ǐ��׏ُ�!�� E�3�i�W���{���ß ���՟����5�G� �g���w�����ѯ�� ����+�=�O��_� a�s�����Ϳ߿�� ��'��K�9�[�]�o� �ϓ��Ϸ�������� !�G�5�k�Yߏ�}߳� �����������1�� U�C�y�g���Y��� ������	�+�-�?� u�c������������� ��;)Kq� �O����� 7%GI[� ������/3/ !/W/E/{/i/�/�/�/ �/�/�/�/??A?S? ��k?}?;?9?�?�?�? �?O�?OO+OaOsO �OCO�O�O�O�O�O_ _'_9_�O]_K_�_o_ �_�_�_�_�_�_�_#o o3o5oGo}oko�o�o �o�o�o�o�oC 1gU�y��� �_?��!��Q�?� a���u�����Ϗ��� ��)��M�;�q�_� ������˟������ %��I�7�m�[�}��� ��ǯ���ٯ���� !�3�i�W���{����� տÿ����/��S� A�wω�3��ϳ�9�o� ������=�+�M�s� aߗߩ߻�yߋ����� ��9�K�]�o�)�� ������������ 5�#�Y�G�i���}��� ���������� UCyg���� �������EW /u����� /�)/;/M/_//�/ q/�/�/�/�/�/?? �/7?%?[?I??m?�? �?�?�?�?�?�?!OO EO3OUO{OiO�O�O�O �O�O�O�O�O_A_/_ e_S_�_w_�_�_i�_ �_�_�_+ooOo=o_o aoso�o�o�o�o�o��o'K9oY~ s �p�s �v���r�$TBJO�P_GRP 2"�au� / ?��v	�r�s�$�|�ip��@� �0�u  � �� � � �=�t @�p�r	 �BL  I�?Cр D�w�q�e�>�n�j�|�<��B$?����@���?�33C�S���a���ǇI�[�x}����;�2�������@��?���z;���V�A�g��〝 ���6�ƕp>̧�����;���pA:�?�ff�@&ff?�ff��ޟa� ��u�󄦁x��,�:v,���c?L����ʐDH�x^�d�v�@�33�����>ʐ������8���퉡�q=�2�D"�����������x=�9�K�9��ݯ ﯐�������חɿ�� ��� �����?�Y�C� Q�ϰϋ�E�������0���@ߙsC��v2����	V3.0~�	lr2d�t�*���t�q�ߤ�� E8� EJ�� E\� En�@ E�pE�� �E�� E�� �E�� E�h �E�H E�0 �E� Eϻ���� E��� �E�x E�X �F���D�  �D�` E���P E��$��0���;��G��R��^op Ek��u�����І��(��� �E��Н�УX O9�IR]�)�q��������v���9�՟���tESTPARSr��x�p�s�HR��ABLE �1%�ys��tD��� `��������w�q��	��
�����.��q�������t��RDI��q-�?�Q�c�u�����O��	%7HI[�S���s �� .@Rdv�� �����//*/ </N/`/r/�}� ��r ,��)����~�������������"NUoM  au�q%��p s�t��_CFG &�;�/3=�@�pIMEBF_TT��*5�s���6VERr��!�6��3R 1'� �8�ߙr�p7A dp�/  O1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_�_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[���� �����!�3���RA_|1�6@�5��MI_CHAN�7� �5 ��DBGL�Vڀ�5�5�ᡀE�THERAD ?U������G��E����血ROUmT�0!�
!S��q�D�SNMASK���3��255.���wӭ���џw���O�OLOFS_DI���k�ӉORQC?TRL (Kg��O�T>�s������� ��ͯ߯���'�9� K�]�o�������=�ƿ������PE_DE�TAIǈ�PGL�_CONFIG �.�9�1��/�cell/$CID$/grp1�@d�vψϚϬ�b�:� ��������1���U� g�yߋߝ߯�>����� ��	��-����c�u� �����L������ �)�;���_�q����� ����H�Z���%7I�.}��������G1ۿ�� ��6HZl~��� �����/�2/ D/V/h/z/�/�/-/�/ �/�/�/
??�/@?R? d?v?�?�?)?�?�?�? �?OO*O�?NO`OrO �O�O�O7O�O�O�O_ _&_�OJ_\_n_�_�_ �_�_E_�_�_�_o"o 4o�_Xojo|o�o�o�o Ao�o�o�o0B�=��User� View R�}�}1234567890s����`��t^�2����Yy2fy�o7�I�[�m������`r3�ߏ���'�9���Z��4 Ώ������ɟ۟�L���5��G�Y�k�}� ���� �¯�66��� ��1�C�U���v��7꯯���ӿ���	�h�*��8��c�uχ���ϫϽ������ �lCameradzZ�#�5�G�Y�k�}�[Eߧ߹��� q����	��-�?�5�  ���ߏ��� ���������1�|�U�g�y���������� ��͉F���1C U��y������ ��	������� gy����h� �	/T-/?/Q/c/u/ �/.��[� /�/�/�/ ??/?�S?e?w?�/ �?�?�?�?�?�?�/�� 驊??OQOcOuO�O�O @?�O�O�O,O__)_ ;_M___O�����O�_ �_�_�_�_o�O)o;o Mo�_qo�o�o�o�o�o r_��Q�bo);M _qo��������%�7��o�g9 �x���������ҏy ����+�P�b�t�P������9�	��00� ���	��-�?��c� u���.�����ϯ�� ������۩�^�p� ��������_�ܿ� � K�$�6�H�Z�l�~�%� ��r�������� �� $�˿H�Z�l߷ϐߢ� �������ߑ�˕���� 6�H�Z�l�~��7ߴ� ����#���� �2�D� V����J������� �������� 2D�� hz����i�� �+Y 2DVh ������� 
//./��"K�z/ �/�/�/�/�/{�/
? ?g/@?R?d?v?�?�?A-  E)�?�? �?�?O#O5OGOYOkO<}O�K   �?�? �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� ��������L�  
A (  }�0( 	 � G�5�k�Y���}����� Ïŏ׏���1��U�:��J ��/�� ����1?�����*� <�C#��f�x���џ�� ��ү����O�,�>� P���t���������ο ����]�:�L�^� pςϔ�ۿ������� 5��$�6�H�Z�l߳� �ߢߴ����������  �2�y�V�h�z��ߞ� ����������?�Q�.� @�R���v��������� �����_�<N `r������� %&8J\� �������� /"/4/{X/j/|/� �/�/�/�/�/�/A/? 0?B?�/f?x?�?�?�? �???�?OOa?>O PObOtO�O�O�?�O�O �O'O__(_:_L_^_ �O�_�_�_�O�_�_�_� oo$ok_K�@  FbSoeowoFcMg1����+frh:\�tpgl\rob�ots\lrm2�00id�`_ma�te_�b.xml 3o�o�o%7I0[moV���� ������,�>� P�b�t��������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l��� }�����Ưد����  �2�D�V�h��y��� ��¿Կ���
��.� @�R�d�{�uϚϬϾ� ��������*�<�N� `�w�qߖߨߺ����� ����&�8�J�\�n�:�h�Q Mo�`�<< �` ?�n��n�������� �/��G�e�K�]�� ���������������3aoV�$T�PGL_OUTP�UT 1yQyQ/ ���� ����0B Tfx����� ��//,/>/P/�����f 2345678901u/�/�/ �/�/�/�#oRr/�/? "?4?F?X?�/\?�?�?�?�?�?n:}�?OO ,O>OPO�?�?�O�O�O �O�O�OxO�O_(_:_ L_^_�Ol_�_�_�_�_ �_t_�_o$o6oHoZo loozo�o�o�o�o�o �o�o 2DVh  ������� �.�@�R�d�v���� ����Џ�􏌏��*� <�N�`�r�������� ̟ޟ�����8�J� \�n����q}�ᶯ@ȯگ����!�@���E�W��� ( 	 Z/��z�����Կ ¿����
��R�@� v�dϚψϾϬ����� ����<�*�`�N�p�@r߄ߺߨ���h&��� �����*��L�^�8� ���b*������q��� �����C�U���Y��� %�w���������	g� ��?��+u�a� ����); Gq����S ����%/7/�[/ m//Y/�/}/�/�/�/ I/�/!?�/?W?i?C? �?�?�/�?�?�?�?O O�?%OSO�?;O�O�O 5O�O�O�O�O_eOwO =_O_�O[_�___q_�_ �_+_�_o�_�_9oKo %ooo�o�_io�oQo�o �o�o�o#5�ok }�����G Y�1��9�g�A�S� �����ӏ��я�����Q�c���)WGL1.XML!�����$TPOFF_LIM ��+�������N_�SV��  (����P_MON M2��+�+��2��STRTCHOK 3���������VTCOMPA�T՘_�ĖVWVA/R 4����ٔ� 6� ��������_DEFP�ROG %$��%	LABWEL�D_�����_DISPLAY��$�ʢ�INST_MSK�  � �I�NUSERU��L�CK^�%�QUIC�KMEN���SC�RE����`�tpsc�^���h����Ұ_ֹSTS����RACE_CF�G 5�������	��
?��HNL 26٪��A��� ��uχϙϫϽ����������ITE�M 27a� ��%$123456�7890H�Z�  �=<R�xߊߒ�  #!�ߠ۬�\��� ��F��j�*�<��R� ���ߟ��ߺ������ v�f�x����(��� ~��������>�P�b� ����2Xj��v�� ��L� *����� � �6�Z�5/�P/ �`/�/�/��/ /2/ D/�/h/?:?L?�/p? �/�/�/|?�?.?�? O d?O�?�?cO�?~O�? �O�OO�O<ONO_rO 2_�OB_h_�O�O�O_ _&_�_J_�_o.o�_ Ro�_�_�_To�_�o�o �oFo�ojo|o�o` �o���o�0� T�x8�J��`�� $����ȏ,�؏��� t��������6����� ��ğ(��L�^�p��� ���f�x�ܟ�� �� ۯ6���Z��,���B�P��Ư���S'�8-�>���  Ҕ�� 9���
 �����B�úUD�1:\O�����R_GRP 195��� 	 @ 렚Ϭ˖��Ϻ������ޠ$�;�I��O��s�^ߗ߂�?�   ���ۮ��������,� �<�>�P��t������������(�	�b�<�N���SCB ;2:�� �ߚ� ����������*���UTORIAL� ;��6�u��V�_CONFIG <��4��2����OUTPUT y=��� ��� $6HZl~�� ������$/ 6/H/Z/l/~/�/�/�/ �/�/�/�// ?2?D? V?h?z?�?�?�?�?�? �?�?	?O.O@OROdO vO�O�O�O�O�O�O�O _O*_<_N_`_r_�_ �_�_�_�_�_�_o_ &o8oJo\ono�o�o�o �o�o�o�o�oo"4 FXj|���� ����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��� �P�b�t������� ��ο����(�� L�^�pςϔϦϸ��� ���� ��$�5�H�Z� l�~ߐߢߴ������� ��� �2�C�V�h�z� ������������
� �.�?�R�d�v����� ����������* ;�N`r���� ���&8I \n������ ��/"/4/EX/j/ |/�/�/�/�/�/�/�/ ??0?A/T?f?x?�? �?�?�?�?�?�?OO ,O>OO?bOtO�O�O�O �O�O�O�O__(_:_>����Y_k_ UQD_�_9��_�_�_�_ oo&o8oJo\ono�o �oEO�o�o�o�o�o "4FXj|�� �o������0� B�T�f�x�������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϯ� ��������
��.�@� R�d�v߈ߚ߽߬��� ������*�<�N�`� r����������� ��&�8�J�\�n�����������$TX_�SCREEN 1}>mUUP�}�����	-?Q���V���� ����bt!3 EWi{��� ���//�A/� e/w/�/�/�/�/6/H/ �/??+?=?O?�/s? �/�?�?�?�?�?�?h? O�?9OKO]OoO�O�O 
OO�O�O�O�O_#_ �OG_�Ok_}_�_�_�_��_<_�_�$UAL�RM_MSG ?5����� �_�� o-o^oQo�ouo�o�o �o�o�o �o$H~�USEV  
m�zv�RECFG� @���� � ��@�  A��q   Bȶ�
 I������� �%�7�I�[�m��������qGRP 2A�{ 0��	 ����PI_BBL�_NOTE B��zT���l������p��D_EFPRO`%
k (%<c���Q� ��u�����ҟ����ៀ�,��P�;�t��F�KEYDATA �1C��Ӏp �w��֏ٯ�¯��!���,(-�T���(�[ INST �]\�^�  ELDG_ST������P���߿B�CHOICE�w��[EDCMqD��7�B�OREq�FO8�;�xϊ�qϮ� �����������,�>��%�b�I߆ߘ� ���/frh/g�ui/white�home.png�������������inst��R�d�v���)�  ��a?rc_str@�D��������'���weldA�]�o�������>4�choic�������'*���edcmK���hz���/���arwrg@���/ ��L^p���� G�� //$/6/� Z/l/~/�/�/�/C/�/ �/�/? ?2?D?�/h? z?�?�?�?�?Q?�?�? 
OO.O@O�?dOvO�O �O�O�O�O���O�O_  _2_D_V_]Oz_�_�_ �_�_�_c_�_
oo.o @oRo�_do�o�o�o�o �o�oqo*<N `�o������ m��&�8�J�\�n� �������ȏڏ�{� �"�4�F�X�j���|� ����ğ֟������ 0�B�T�f�x������ ��ү������,�>� P�b�t��������ο���ϟ���>�����:�L� ^�6πϒ�l�,~��� v��������A�(� e�w�^ߛ߂߿��߸� �����+��O�6�s� Z���������� �O'�9�K�]�o����� �������������� 5GYk}�� �����1C Ugy��,�� ��	//�?/Q/c/ u/�/�/(/�/�/�/�/ ??)?�/M?_?q?�? �?�?6?�?�?�?OO %O�?IO[OmOO�O�O �ODO�O�O�O_!_3_ �OW_i_{_�_�_�_@_ �_�_�_oo/oAo� eowo�o�o�o�o�_�o �o+=O�os �����\�� �'�9�K��o����� ����ɏۏj����#� 5�G�Y��}������� şןf�����1�C� U�g�����������ӯ �t�	��-�?�Q�c� 򯇿������Ͽ�� ���)�;�M�_�q� � �ϧϹ�������~�߀%�7�I�[�m��V`����V`����߼��ݦ������,��3���W�>�{�� t������������ /�A�(�e�L������� �������� = $asRo���� �� �'9K] o������ ��#/5/G/Y/k/}/ /�/�/�/�/�/�/? �/1?C?U?g?y?�?? �?�?�?�?�?	O�?-O ?OQOcOuO�O�O(O�O �O�O�O__�O;_M_ __q_�_�_$_�_�_�_ �_oo%o�_Io[omo o�o�o2o�o�o�o�o !�oEWi{� �������� /�6S�e�w������� ��N������+�=� ̏a�s���������J� ߟ���'�9�K�ڟ o���������ɯX�� ���#�5�G�֯k�}� ������ſ׿f���� �1�C�U��yϋϝ� ������b���	��-� ?�Q�c��χߙ߽߫� ����p���)�;�M� _��߃�����������p����p����,�>��`�r�L�,^��V�� ��������!EW >{b����� ��/S:w �p�����/ /+/=/O/a/p�/�/ �/�/�/�/�/�/?'? 9?K?]?o?�/�?�?�? �?�?�?|?O#O5OGO YOkO}OO�O�O�O�O �O�O�O_1_C_U_g_ y__�_�_�_�_�_�_ 	o�_-o?oQocouo�o o�o�o�o�o�o�o );M_q��$ �������7� I�[�m���� ���Ǐ ُ����!��E�W� i�{�������ß՟� ����/���S�e�w� ������<�ѯ���� �+���O�a�s����� ����J�߿���'� 9�ȿ]�oρϓϥϷ� F��������#�5�G� ��k�}ߏߡ߳���T� ������1�C���g� y��������b��� 	��-�?�Q���u��� ��������^����);M_6�a}�6�����@������,� �7[mT� x�����/!/ /E/,/i/{/b/�/�/ �/�/�/�/�/??A? S?2�w?�?�?�?�?�? ���?OO+O=OOOaO �?�O�O�O�O�O�OnO __'_9_K_]_�O�_ �_�_�_�_�_�_|_o #o5oGoYoko�_�o�o �o�o�o�oxo1 CUgy��� �����-�?�Q� c�u��������Ϗ� ����)�;�M�_�q� �������˟ݟ�� ��%�7�I�[�m���� h?��ǯٯ����� 3�E�W�i�{�����.� ÿտ����Ϭ�A� S�e�wωϛ�*Ͽ��� ������+ߺ�O�a� s߅ߗߩ�8������� ��'��K�]�o�� ����F�������� #�5���Y�k�}����� ��B�������1 C��gy���� P��	-?� cu����������������/-�@/R/,&,>?�/6?�/�/�/ �/�/?�/%?7??[? B??�?x?�?�?�?�? �?O�?3OOWOiOPO �OtO�O�O���O�O_ _/_A_Pe_w_�_�_ �_�_�_`_�_oo+o =oOo�_so�o�o�o�o �o\o�o'9K ]�o������ j��#�5�G�Y�� }�������ŏ׏�x� ��1�C�U�g����� ������ӟ�t�	�� -�?�Q�c�u������ ��ϯ�󯂯�)�;� M�_�q� �������˿ ݿ���O%�7�I�[� m�φ��ϵ������� ��ߞ�3�E�W�i�{� ��߱���������� ��/�A�S�e�w��� *������������ =�O�a�s�����&��� ������'��K ]o���4�� ��#�GYk }���B��� //1/�U/g/y/�/ �/�/>/�/�/�/	??h-???�A;�����j?|?�=f?�?�?�6,�O�?�O O�?;OMO4OqOXO�O �O�O�O�O�O_�O%_ _I_[_B__f_�_�_ �_�_�_�_�_!o3o� Woio{o�o�o�o�/�o �o�o/A�oe w����N�� ��+�=��a�s��� ������͏\���� '�9�K�ڏo������� ��ɟX�����#�5� G�Y��}�������ů ׯf�����1�C�U� �y���������ӿ� t�	��-�?�Q�c�� �ϙϫϽ�����p�� �)�;�M�_�q�Ho�� �߹����������%� 7�I�[�m����� ���������!�3�E� W�i�{�
��������� ������/ASe w������ �+=Oas� �&����// �9/K/]/o/�/�/"/ �/�/�/�/�/?#?�/ G?Y?k?}?�?�?0?�? �?�?�?OO�?COUO@gOyO�O�O�O���K���������O�O�M�O _2_V, oc_o�_n_�_�_�_ �_�_oo�_;o"o_o qoXo�o|o�o�o�o�o �o�o7I0mT ��������� !�0OE�W�i�{����� ��@�Տ�����/� ��S�e�w�������<� џ�����+�=�̟ a�s���������J�߯ ���'�9�ȯ]�o� ��������ɿX���� �#�5�G�ֿk�}Ϗ� �ϳ���T������� 1�C�U���yߋߝ߯� ����b���	��-�?� Q���u������� ����)�;�M�_� f�������������� ~�%7I[m�� ������z !3EWi{
� ������/// A/S/e/w//�/�/�/ �/�/�/?�/+?=?O? a?s?�??�?�?�?�? �?O�?'O9OKO]OoO �O�O"O�O�O�O�O�O _�O5_G_Y_k_}_�_ _�_�_�_�_�_oo���!k������Jo\onmFo�o�o|f,��o��o�o -Q8u�n �������)� ;�"�_�F���j����� ��ݏď����7�I� [�m�����_��ǟٟ ����!���E�W�i� {�����.�ïկ��� ����A�S�e�w��� ����<�ѿ����� +Ϻ�O�a�sυϗϩ� 8���������'�9� ��]�o߁ߓߥ߷�F� �������#�5���Y� k�}������T��� ����1�C���g�y� ��������P�����	 -?Q(�u�� ������) ;M_����� ��l//%/7/I/ [/�/�/�/�/�/�/ �/z/?!?3?E?W?i? �/�?�?�?�?�?�?v? OO/OAOSOeOwOO �O�O�O�O�O�O�O_ +_=_O_a_s__�_�_ �_�_�_�_o�_'o9o Ko]ooo�oo�o�o�o �o�o�o�o#5GY�k}��$UI_�INUSER  �����q�  ���_MENHIS�T 1D�u�  ( ��p��./SOF�TPART/GE�NLINK?cu�rrent=ed�itpage,L�ABWELD_2�,1�H�Z�l�z)�	��menu'�16315�ŏ׏���' �'����7��F��X�j�|�r(���95,18��Ο���������,148,2�R�d�v����)�,1546�ԯ����
�p/���AB_ /�5�^�p����#�5��G�4�������� p�(�3�E�W�i�{��ϟ� /��������� �߭�B�T�f�xߊ� ��+����������� ,��P�b�t���� 9���������(��� L�^�p���������G� ���� $6!�Z l~������� � 2D�hz ����Q��
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?�/r?�?�?�?�? �?�?m?OO&O8OJO \OGeO�O�O�O�O�O �O�?_"_4_F_X_j_ �O�_�_�_�_�_�_w_ �_o0oBoTofoxoo �o�o�o�o�o�o�o ,>Pbt�� ������(�:� L�^�p���mO���ʏ ܏� ���6�H�Z� l�~������Ɵ؟� ��� ���D�V�h�z� ����-�¯ԯ���
� ���@�R�d�v����� ��;�п�����*� ��N�`�rτϖϨϓ���$UI_PAN�EDATA 1F�������  	�}�/frh/gui���dev0.st�m ?_widt�h=0&_hei?ght=10	����ice=TP&_�lines=15�&_column�s=4	�font�=24&_page=whole����ϑ�)primX߁�  }�ߨߺ�0������� )�(� �L�3�p��i��� ������ ���$�6���Z����� �  z��" �ߗ�����������D� ��9K]o�� �������# 
G.k}d�� ����n� ��% ��6;/M/_/q/�/�/ ��/,�/�/??%? 7?�/[?m?T?�?x?�? �?�?�?�?O�?3OEO ,OiOPO�O�O/$/�O �O�O__/_�OS_�/ w_�_�_�_�_�_�_J_ o�_+ooOoaoHo�o lo�o�o�o�o�o �o9�O�Oo��� ����r_#�5� G�Y�k�}������ŏ ׏������1��U� <�y���r�����ӟF X��-�?�Q�c�u� ȟ�����ϯ��� �~�;�M�4�q�X��� ����˿���ֿ�%� �I�0�m������ ���������b�3ߦ� W�i�{ߍߟ߱���*� �������/�A�(�e� L���������� ����Ϟ�O�a�s��� ����������R� '9K]���h� ������5 YkR�v�&�8�}���/!/3/E/W/)�|/��k/�/ �/�/�/�/?i/&?? J?1?C?�?g?�?�?�? �?�?�?�?"O4OOXO���B�<��$UI_�POSTYPE � B��� 	 dO�O�BQ�UICKMEN � �K�O�O�@R�ESTORE 1�GB�  O�KO��5_BS0_��m`_�_�_�_ �_�_t_�_oo+o=o �_aoso�o�o�oT_�o �o�oLo'9K]  ������~ ��#�5�G��oT�f� x����ŏ׏����� �1�C�U�g�
����� ����ӟ~�����v� (�Q�c�u�����<��� ϯ�����)�;�M� _�q��~������ݿ ���%�ȿI�[�m� ϑϣ�F��������ϼ��GSCRE�@?��Mu1s]c*Pu2J�3J�U4J�5J�6J�7JԹ8J�'�TAT�M�� �CB��JUSE�R,�1�C�T+�L�k�sT���4��5��6���7��8�ъ@ND�O_CFG H��K���@PD������Non�e�B��_INFOW 1IB�q��@0%ߌ���z��� �������'�
�K�.� o���d����������L�^�OFFSET L�Iu�����#P ��,>Pb��� ����( UL^������O��/
/:/���UFRAME  ���.�[�RTO?L_ABRT^/Y��v"ENB/p(GR�P 1MY�ACz  A��#�!3� �/�/�/	??-???Q;�r&�@U�(3�+MS�K  �%q�+N6[!%i��%��?��%_EVN~ �4�-��6�2N

 }h3�UEV~ �!td:\ev�ent_user\�?B@C7GO/��YF|L:ASP@AEG�spotweldwM!C6�O}O�O*P�4!�?VO_I_�G �1_8_&_|_�_\_n_ �_�_o�_�_�_So�_ wo"o4ojo�o�o�o�o �o�o+O�o� 0��fx������zFWRK 2O��&!8�y��� g��������ӏ �.�	�R�d�?����� u���П������*��<��M�r����$V�ARS_CONFuI"�P
 FP�û���CMR�"2�V
�9��	�4ೠ��1: S�C130EF2 Q*���ę���x֊0�5��3�?��a0@a0pU0ȅ� )/h�r��ȓ�@��ҿ��Ϳ��k�O5�A���7ϲ�? B���R��� V�޿wϾ���jϿϪ� ��������=ߔ�� s�^�pߩ�\����ߓ��IA_WOQ�W<i��v,		�F�|(�6�G�P �I���H��RTWINU_RL ?&I����ߎ������������SIONTM;OUO � �B�XS۳�S���@�! FR�:\�\DATA��O  �� �MCA�LOGN� �  UD1A�E�Xr���' B@ �����`�����������x �� n6  �������6��  =���M�J ���g�TRAINМ�\�Bd�p�MQ����ңY&K (�ѝ	����� %[Im���������_GuE)�Z&K�`
���
� 
�?"'��R�E,�[�)����LE�X $\���1-e���VMPHASE'  &E�N����RTD_FILT�ER 2]&K �1��_� ??$?6? H?Z?l?~?�?�?��/ �?�?�?OO*O<ONO�`OrO��SHIFTMENU 1^�/
 <��%���O����O�O_�O�O C__,_y_P_b_�_�_��_�_�_�_�_-oo�	LIVE/SN�A��%vsflsiv�.?o�� SETU��bbmenuxo}oo�o�o�#�E)�_k�HMO�)�`.�z��ZD�ta\/
�<��P��$WAITDINEND��!rvvOK  ꩑|�r�S��yTIM����|G}���0�������xRELE�!@�vvs�<�xq_ACTU`?�t�x_J� b���%�o@����RD�IS����vpV_oAXSR|�2cYy�w�D(|�Ӡ_IR 3 �&t� 7
ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚϸ�Ͼ�NXVRy!�d7~�$ZABCv�1eY{ ,� �2����Oq��VSPT f7}�r{�
�j�o���j��ߣ�B�DCSCHb{ g�d���IPRrhY�6�H�Z��l���MPCF_G 1i��05׫�q�MP�j�6 �p5�����<��0  ?t�?/��>�����*?����Mو�I��R>�ԅ>��}C��CB�_�Õ���?��@�?������I�?�Bc��� ����$�6�H�1V�h�z����������/��� �D�B��jA{"�v�2���EC
#�FX?����������~�O��'}&&�y�3\�L��3���Q?���.��C�����_5�$����0.� �ڽ�Z��{ �k�W_CYLI�ND�!l�� ���� ,(  * ���Ӧ��/� 4=/O/a.��/ ��/�/�/�/!/?? &?i/J?�/�/�?g?�?��?�/�?�?O��2md� ġ�7OGL j�3pO[O�O��'O�Oʹז�AA��ySPHERE 2n��>?_�?_P_7_t_ �?�O�_�_8?�__e_ o�_:o!o�_po�o�_ �_�o+o�o�o�oYo�6HZ��ZZކ �ʆ