��   ��A��*SYST�EM*��V9.1�0214 8/�21/2020 A 
  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41�� d =R��&J_�  4 $:(F3IDX���_ICIgMI/X_BG-y
�_NAMc MO�Dc_USd�I�FY_TI� �MKR- � $LINc  � "_SIZ��$�� �. �X $USE_FLC 3!�:&iF*SIMA7#QC#zQBn'SCAN�[AX�+IN�*I���_COUNrRO�( ��!_TMR_cVA�g#h >�ia �'` ��p��1�+WAR�K$�H�!�#N33CH�PE�$O��!PR�'Ioq6��OoATH- �P $ENABL+�0BT�ELD�$$CL�ASS  �S���1��5��5�0�VERS��7  �AIRTU� �?@'|/ 0E5���E����@kF1@�1pE��%�1�O���O��O����AEI2LK�_,_>_P_b_ t_�_�_�_�_�_�_�_�oo(o:o�O*W?yHW@ �� zj�0�o�o�i�� �� 2LI  #4%Ho�o��mA}A �o+
Oa@��v���@�A��� �(���^�=�1@�c�$"+ �k�K@����pA��XmA0A@ �N�����0�B�T� f�x�����������pF }AՁ}A����*�<� N�`�r���������̯�ޯ�4hL��C� 2�lՏ;�M� _�q���������˿ݿ ���Ԝ-�F�X�j� |ώϠϲ��������� ��)�B�T�f�xߊ� �߮����������� ,�7�P�b�t���� ����������(�3� E�^�p����������� ���� $6A�Z l~������ � 2DOhz �������
/ /./@/K]v/�/�/ �/�/�/�/�/??*? <?N?Qh�4�0���?�p