��   g�A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG  �DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST� �DwNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !���FT�{ @� LOG_8	�,CMO>$D�NLD_FILT�ER�SUBDI/RCAPC � �\8 . 4� H�{ADDRTYPz�H NGTH�̉��z +LS�q D $R�OBOTIG �P�EER�� MAS�K�MRU~OM�GDEV����P�INFO� � $$$TI� ��RCM�+T A$x( /�QSIZ��!S� TATUS�_%$MAILS�ERV $PL�AN� <$LI}N<$CLU��ި<$TO�P$�CC�&FR�&YJ�EC|!Z%ENB{ � ALAR:!�B�TP,�#,V�8 S��$VAR�)M�ON�&���&oAPPL�&PA� 8�%��'POR�Y#�_�!�"ALERT��&i2URL }}Z3ATTAC���0ERR_THROU3US�9H!�8� �CH- c%�4MAX�?WS_|1�N�1MOD��1I� � �1o (�1PW7D  � LA��0v�ND�1TRYFDELA-C�0G'A�ERSI��1Q'R]OBICLK_HM 0�Q'� XML+ 3S/GFRMU3T� !3OUU3 G_�-C�OP1�F33�AQ'C8[2�%�B_AU�� p9 R�!UPDb&�PCOU{!�CFO� 2 
$Vp*W�@c%ACC_H�YQSNA�UMM�Y1oW2��RD�M*� $DI�S��SM	C l5�o!�"%Q7��IZP�%� �VR�0�UP� _DLV�SPAR�SN,#
3 �_�R!�_WI�CTZ_I�NDE�3^`OFF,� ~URmiD�)c��   t 9Z!`MON��c�D��bHOUU#E�%A�f�a�f�a�fLOsCA� #$NS0oH_HE���@�I�/  d8`A�RPH&�_IPFF�W_* O�F``�QFAsD90�VHcO_� 5R42PSWq�?�TEL� �P���90W�ORAXQE� L�V�[R2�IC�E��p� �$cs ? ����q��%
��
�p�PS�A�w�  �5�	�Iz0AL��X' �
���F�����!�p�i��$.� 2Q� "���������� Q���!��q����$� _F�LTR  �\�� �����������$Q�2��7rS�H`D 1Q�" P㏙�f���ş ��韬��П1���=� �f���N���r�ӯ�� �����ޯ�Q��u� 8���\�������󿶿 �ڿ;���_�"�Xϕ� �Ϲ�|��Ϡ����� ��6�[���Bߣ�f� �ߊ��߮���!���E� �i�,��P�b���� ������/���(�e��T���L�����z _L�UA1�x!1E.��0��p���1��>p�255.0��&r��n���2����@d %7I[3e���� ����[4 ���T'9[5U���{���[6���D �//�)/s��QȁM�A¸MA�H������ 'Q� ��u.<�/? &?�/J?\?n?A?�?�?m�P�?�?�?�?�?O .O@OROOvO�O�Ou.�kOl�q��O�L
�ZDT StatusZO�O5_G_Y_n��}iRConn�ect: irc�{T//alert ^�_�_�_�_mW#_o@o,o>oPobot�^�P~2g���go�o�o �o�o�o�o	-?�Qcul�$$c9�62b37a-1�ac0-eb2a�-f1c7-8c�6eb5189a8c  (�_�_ ���"�p�1!W��(��"S��JE�� 0X��C� ��,$��� W���ˏ���֏�� %��I�0�m��f��� ��ǟ�������!���u�R����� D�M_�!����S�MTP_CTRLg 	����%� ���DF���ۯt�ʯ���'��Lz�N��!
�j��y�q�u�����Ԙ��#L�US?TOM j�������  ���$T�CPIPd�j���H�%�"�EL������!���H!T��b<�n�rj3/_tpd7� ��i�?!KCLG�L��i���5�!CRT�ϔ����"u�!OCONS��M�[�ib_smon����