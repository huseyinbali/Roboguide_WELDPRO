��   v��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@ � &�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	�c&USRVI| 1  < `��R*�R��QPRIƍm� t1�PTR�IP�"m�$$C�LASP ��)�a��R��R `\ �SI�	g�  �aIR�Ts1	o`'2 L1���L1���R	 �,��?����a1`�b�d~a����c��y`� � ����
 ���'/SOFTP��@/GEN�1?CURRENT=>>�A,18,1�o�1CU �o�o,95,2W����' �(k}5	p��(�:�L�^�i��q9 _�����Ϗ������/�A�S�e���E,381��ğ֟ �o�a��%�7�I� [�m���������ǯٯ �z��!�3�E�W�i� ��������ÿտ����~aTPTX������/�` �sȄ�$/so�ftpart/g�enlink?h�elp=/md/�tpmenu.dg���ϨϺ��υ��� ��&�8�J���n߀� �ߤ߶���W������ "�4�F�X���|��ﰲ��������a�f�b�b�� ($ p�-����T�?�x���a�a��c���g��Il��k
��ah�*�ah�h�2�h�]	f����������`���`  ����f epT��h#h�Fd��g��Xc�B 1)hR� \ _�b� REG V�ED]���wh�olemod.h�tm�	singl�	doub �trip8browsQ�� ���u���/�/@/���dev.sl�/3� 1�,	t�/_�/;/ i/??/?�/S?e?w?8�?�?�?� H`�? �? OO$O6OHOZOlO ~O�F2P�?�O�O�O�O �O_�E�	�?�?;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo oM'�o�o�o�o�o�o +=Oas� ��������? >�P�b�t��������� Ώ���O�����L� ^�_'_�������ş �����6�1�C�U� ~�y�����Ư��ӯ�o ���-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�-��Ϭ� ����������*�<� 7�`�r�A�Sߨߺ�q� ��i�����!�J�E� W�i��������� ����"��/���O�I� w��������������� +=Oas� ������, >Pbt���߼ ���//����� ^/Y/k/}/�/�/�/�/ �/�/�/?6?1?C?U? ~?y?�?Y��?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _�R_d_v_�_�_�_ �_�_�_�_�o*o�_�o`oro�j�$UI�_TOPMENU� 1K`�aR 
d�a�*Q)*defa�ult5_]*�level0 * [	 �o�0��o'rtpio�[23]�8tpst[1[x)w9��o	�=h58E�01_l.png���6menu5�y�p�13�z��zb	�4���q��]� ��������̏ޏ)Rr����+�=�O�a����prim=�pa�ge,1422,1h�����şן����1�C�U�g����|�class,5�p�����ɯۯ�����13��*�<�N�`�4r���|�53�������ҿ�����|�8 ��1�C�U�g�y�����@����������"Y�` �a�o/��m!ηq�Y��w�avtyl}Tfqm�f[0nl�	��c�[164[w��59@[x�qG���/��29� �o�%�1���{��m� �!�����0�B��� f�x���������O������,>����2 P�����\�� '9K�������������1���/$/6/H/Z/��~|�ainedi'���/�/�/�/�/��c�onfig=si�ngle&|�wintp���/$?6?H? Z?!Z�a�h?�?�e�? �;��?�?�?OO+O =OOO�?[O�O�O�O�O �O�O�O_a�%_L_^_ p_�_�_�_���_�_�_  oo$o�_HoZolo~o �o�o1o�o�o�o�o  2�oVhz�� �?���
��.� �@�d�v��������� M�����*�<�ˏ�`�r���������^ ��;�M�sc�_;����s��X�}���e�u ��0���P��t���4�j�X�6e�u7 �����ｿϿ��� P�)�;�M�_�qσ�� �Ϲ����������"�1�M�_�q߃� �ߠϹ��������� ��7�I�[�m���� ����������!�����6(�]�o��������$��74�������)t<ϯ\�5	TPTX[209©|Dw24§J����w18����
�02��A#��[�tv`�RdvL0�K1���5S�:�$treevi�ew3��3��&d�ual=o'81,26,4�O/a/ s/2�/�/�/�/�/�/ �/?'?9?K?]?o?��;/��53$/6$�� �?�?�?
?#O5OGOYO kO}OO�O�O�O�O�O��O�?�?��1�?6$2p�f_x_�_ �6_��edit��>_P_ �_�_o��/���_�S ooo�o�oB�o�o� �oA�o�+= Oas��o��� ����(�9���Q� x���������ҏ�O�� ��,�>�P�ߏt��� ������Ο]����� (�:�L�^�ퟂ����� ��ʯܯk� ��$�6� H�Z��l�������ƿ ؿ�y�� �2�D�V� h����Ϟϰ������� �o�o��o@ߧE�c� u߇ߙ߽߬�����O� ���)�<�M�_�q�� ��W���������&� 8���\�n��������� E�������"4�� Xj|����S ��0B�f x����O�� //,/>/P/�t/�/ �/�/�/�/]/�/?? (?:?L?��߂?1ߦ? ���?�?�?�?O$O 5OGO�?SO}O�O�O�O �O�O�O�O��2_D_V_ h_z_�_�_�/�_�_�_ �_
oo�_@oRodovo �o�o)o�o�o�o�o *�oN`r�� �7�����&� �J�\�n��������� E�ڏ����"�4�Ï X�j�|�������a?s? 蟗?�sO_/�A�S� e�w����������� ����,�=�O�a�#_ ������ο��=�� (�:�L�^�pς�Ϧ� �������� ߏ�$�6� H�Z�l�~�ߐߴ��� ��������2�D�V� h�z���������� ��
����@�R�d�v� ����)����������ƚԔ*def�ault%��*?level8�ٯ�w���? t?pst[1]�	��y�tpio[#23���u����J\menu7_l.png_M|13��5�h{�y4�u6� ��//'/9/K/]/�� �/�/�/�/�/�/j/�/�?#?5?G?Y?k?�"�prim=|page,74,1p?@�?�?�?�?�?�"�6�class,13 �?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo�]ooo�o`�$UI�_USERVIE�W 1֑֑�R 
��EDIT,We�ld DATA ���double�����obmedit�1�o0BT�j�695�Pa� ���m ��$��6����cSTATU�S,POS�ftrip�o�o�o����ʏ(܏��y2��+�0=�O�a��33�_�� ����ϟz�ܟ� ��� �E�W�i�{���0��� ïկ������/�A� S�e��r������ѿ ����ϼ�=�O�a� sυϗ�:ϻ������� ߮��"�4ߦ�o߁� �ߥ߷�Z�������� #���G�Y�k�}��:� D����2�����1� C�U���y��������� d�����	-��: L^������� �);M_ �����v�� �n7/I/[/m//"/ �/�/�/�/�/�/?!? 3?E?W?/?v?�?�/ �?�?�?�?OO�?AO SOeOwO�O,O�O�O�O �O�O�?__&_�Oa_ s_�_�_�_L_�_�_�_ oo'o�_Ko]ooo�o �o6b