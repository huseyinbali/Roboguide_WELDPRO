��  	G��A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �me�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@  �ALRM�_RECO" � � ALM�"EN5B���&ON�!� �MDG/ 0 �$DEBUG1PA�"d�$3AO� �."��!_IF�� � 
$ENA�BL@C#� P djC#U5K�!MA�hB �"�
� OG�|f 0CURR_D1:P $Q3LIN@S1�I4$C$AUSOd��APPINFO;EQ/ �L �A ?1�5/ �H �79EQUIP 2�0�NAM� ��2_�OVR�$VE�RSI� ��PC�OUPLE,  � $�!PPV1C#ES C G1�2�!�PR0�2	 � �$SOFT�T�_IDBTOTA/L_EQ� Q1]@�NO`BU SPI_OINDE]uEXBSCREEN_�4�BSIG�0�O%KW@PK_FI�0	$THK�Y�GPANEhD �� DUMMY1"d�D�!U4 Q!�RG1R�
 � _$TIT1d  ��� 7Td7T� 7TP�7T55V65V75V8
5V95W05W>W�A7UPRWQ7UfW1pW1zW�1�W1�W 6P����ASBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"=$Nb_OPT�2� �� ELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1�0UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t�
��WELDH2/0 =s�q"Q7ING�0$�QAx7PD2�4%$ASd3��BEl�P�_��BU�CC_AS�BFA�IL��DSB��F3AL0��ABN@��NRDY���`��zv��YN��SCH���pDE���yp���p�����|�STK>�0��	���	�NOj�?�ڂL��d�U* G��� 9 ���������߇ƗpƗ��ԘS_Fә1E��F�ƗSSŘ���P�1 �ON�F�HkOU�D�MI�1D�SEC`B�yi �HEK0~��GGAP������I� Ν GTH���0D_ȡ����T= ��륌� 
��p}�9!K���9!ƗUN14��5��#�MO� �sE �� [M�s��t�R�EV�B�����!X�I� g�R  �� OD}`��ii�`M�a����/�"��� �ŵ�eaX�@Dd� p E RD_�E���$FSSYB�&W`KB!�E2u#AG� J��  "��S�� V�t:5`�QC�`�a_EDu �� � C2�f�S�pa�l �t$OP�@QB�q��_OK<"�آTP_C� ��p�da�U �`LACm��^��J�� FqCOM	M� K�D��р@�p���OR�BIGA�LLOW� (tK\��@VARw�xd!�A}!�BL[@S � ,KJq��rH`S�pZ@M_O]��՗�CFd X�0GR@��=M�NFLI��ӂ;@Uɠ�84�"� S�WI�&"AX_N�o`����9��G�� �0WARNMxp�d4�%`L�Tb;��� COR-rF�LTRY�TRAT� T�`� $AC�C@�TB� ��r�$ORI�.&�R�T�`_SFg� C�HGV0I���T���PA�I��T��e`5��� � ��#@a"��HDRՃ7�2�BJ; �CO�I�3J�4J�5J�6*J�7J�8J�9��Ȱ�x@�2 @� TRQ��$%f�������_U������Oc <� �����
�3�2��LLEC���o�MULTI`V4�"fѱA
2FS�GILD��
1;�Oz@�T_1b  4� STY2�bv�=��)2_��:��� |9$�.pڰ�x�I`�* �TOtF �sE�	EXT�3ء�B3�22X�0��@�	01b.'.�Bp�
���  �"��/%�a@�g�?s��!��;AآM�`Q�  �TRE� " L�0�	�`���pA�$JOB`��E����$IG� # d�,/>/P(����#��_M�ORc$ t�F�͠�CNG�AŠTBA �6c�:/�9@��0�19@G;P/pXH5��?�%L�����Bq�1��&rJ��_!R������;J@��8
�<J� D81��9Q��2�@��;�Rd&� 
	�r�G�R�`HANC?$LGw��a2q� ͠�Z�/��
0�2�R��Li��D��)�f�CDB`�CRA�c�CAZ�`�HELT���FCT<�".�F"�`�M#@�AI([O(X����
1@�Rw�w 3/�S���1��5�MP������HK&AES_S�H�Q�W��N0S���Z����'  �v@I#�Aq�Rc(>��STD_C�t�Q��3"UST�U:��)kTIT�a~�ڤ	%�1IOy����@_Up�q��* \����UpORzs`b���}�~p�`O~@N�SYR�G`�q�eUp�а��� ��G`P_XWORK��+r �$SK��<�p1D�B�TR�p , ��0A���c�B��fW�DJDS _Cd�0`�sDPwPLzq�ё�s��DM�<wY�!���2��H�9N�p�# Eb�A��-�bHa�PRi�M�

�D8�� ��. q��1�$�$Z���eL�y/������r��0����P�� 1��tENE��� 2���a���v��r3H {$C��.$L`��/$�s���tw�IN�EV�a_D}�m�RO3���I;�~!�`��:���RETUR�N���MMRj"U�琋�CʠNEWM�A`#�SIGN��A�J@#�LA<�!�&P�0$Po 1$�P�@�24�M� ;�O��S���a�o���v�Q�V�GO_AW�T #�`�@`ъQWg�DC)�o�CY� 	4'"�1�(����Ĕ2��2̖Na���C��4��DEVI�� 5 P $��RBU��PI̗P<��3�I_BY�;��J�T�1�HNDG�q6 Hv�c&�E�g㸣�#�㗣͖h�`���L�7w���`�Ѭ�FBڬ(�FE�����͔��@�ܱ�8� �МQ��@�MCS4�Ƞ�dH����RHPWF��5:�J �n���SLAV.�9�INP��J���������:P +B�S6@`�� B�� ,1�FI(b�� 	��5OaQ'OaW	�'NTV�V��7SKI�CTE*�@�0��b�]�QJ_S�R9_���SAFv�5���_SV2EXCSLUv`-�D~`�L���Y�{�H�I_VRP�RPPL�Y4px���u�۶��_�ML�v`$VR�FY_s��M�I3OC\�%C_>PS�dT�]�O/���LSр���nt4Fqy�͓�� �`P�en⯐K�AUNF����͕��8�ZqCHD�$������� AF� CPU#��TFqĳ?Pס' ;4��`T��c.�� ��N��' <��8@TЀ��q ��g�óSGN=�0
$U0����� �Б� *0e �b��b>��ANNUN��� ��͕U0�4v`'�w �����>P�����EF�`I�>��$F��&dO0OT��nt@��prTq��kq)�M��NI�r?'"|�G~�Aޱ��DAYecL�OAD�ctu�os5�v�EFF_AXIJɢ@4�Yq�SO��|�s�`_RTRQ�GA Dy�Q� Qt` E����� @�P�WP  ���AMPC@E�� B�XT]2Xl��8FDU�8E��bC�AB�C8�*�NSlj0ID�!WRBhU�A:PV%�V_T � �@�DI%0cD�� 1$V�SE�T�2]3�1�o�0
��]2�1E_��l�VEP	0SW�AQ�0� 3  A�N0��OHqPPLAmIRAa]2B�` �n�����S���@�@�%�� C��P ��RQDWf�MS�P%AXt</lLIFEp�. uq:"NA!M2J%��?#M2C����C�P���N�$ǁ�&��O�V��V&HE��]2S�UP�!��:"p_�$��y!_:3�%���'Z�*W�*�Q�'S�ገ��RXZ�@�qY2=8C��T�`��	QN?���J%Q �a_�@j�� CT�T�E `�CACqHt��3SIZp&� ��%�NZ�UFFI� �p��ct$��os6wry�M�P%D�F 8��KEYI7MAG�TM���C�#A��F��Ɓx�OC'VIEK�aG�R�@�LCĐ� �?� 	R#�D?P�4H b�STo�!�B�ГD�Tp�D��D��@EMAIL�𽀣����/FAUL�rI�R���cPCOU�PFA�`�TO��QJ< �$�C5�ST � IT��BUF�7 ��7
��4`*`� B*T5�C������BAcPSAV uU7R \2:�U�W�����P|T5�R�L��_0*P[U���YOT���`���P2�\p�Z?��WAXec+�=�X*P�éS�_GA#
� YN_\���K <� D0�T!p���M�� 5T��Fƀ$݀��DI �E�`O�P��aIL����GKQF�&������a������	�Ma�\��a�C�SC_���K���`���d��RpA�e�H�aDSP3F6�bPC*{IM�S!sGq��a� U�g� ��"��@IPD��c{0� tTH[0��r��T̩�!sHS�csBSCQ�j0*�Vְ�z�p�!c�tf���NV��G  ��t[0v*PFAB`ads}`aǁSC��&��cMER��bqF�BCMP���`ETn�� NBFU� �DUP���22��CaDy�p�P�CG�ЀSNO�х�O ������PN�C"j�υR�@b�A��|�P��PH *ρL۰����QL���� o�B���@�j�@���@�P��@��1@�7=�8=��9=�A ?�I�1V�1�c�1p�1}�1��1���1��1��2��2TI�V�2c�2p�2}�U2��2��2��2���3��3I�3V�c�3�p�3}�3��3��3ʤ�3��4��DaEX	T���QTb��Y`m&�Y`:�d`����AFD�R�RT
PV����R:"ɱ�r:"RE�M#FU�OVM��c�A��TROVf��DT�P�MX'��IN��� ��IN	D6�
bȎ`B`W`�G*a�!��@J%0D!�RIV�n"oGEAR�aIO'	K�lN}`����%(�L�?@� mZ_MC�M50:!�F� U�R{�S ,́MQ?g � \p?4�.@?4�Et�<�"��gQX���T�0�5Pa� RI�����7SETUP2_ gU ��6STD�px5TT��LѢל��A�7RBACNbV T(��7R�d)�j%<��x`�IFI�x`X��)�A ��PTM��L{UI~DW �� `H PUR�`Q�"�R��a�p-P�$ Iܴ$�p�S$�?x|�J�`CO�P�SVRT|l�G�x$SHO#���CASS�p�Qp%�p��BG_���V����c���p���}�FO�RC�B-�DAT�A��X�BFU�1��b"�2�a*�[0��Y� |r�NAV`S�p����S�B~n#$VISI��6vbSCdSEZм�V��O���B��I� ��$PO�t�I��FM�R2��Z  Ȳ���ɱ�`��ͷ��@������@�_��9��$IT_ᛄ�"M�Ʋ���DGC{LF�DGDY�LDLѐ�5R&��J$R��M���C[G@;	? T�FS�PD�\ Pz��cB`�$EX_.1P`��"3P5Ps�G�q��] �L��x�SW^UO�DE�BUG���GRt��4@U?�BKUJ��O1� O P�O ��j���Mλ�LOOc�SM�K E�R�AT�� _E� ^ 7@��_�TERM %_)%���ORI�ar% `)%�ASM_�`���% a)%��h(b�B&�0UPUBc�3 -S��^p�7#ʮ _��G�*� EL�TO�A�b�FIG�2�aЛ,@N$�$�`$UFR�b�$À�!0��V OT�7�TA�pɰ13N;ST�`PAT�q�0�G2PTHJn���Ep�@�R���"ART�P��%�@�Q�B�aREL<�:9aSHFT�r�aM1{8_��Rw���f&% q $�'�0bvʰ8��\s9bSHI�0s�U9� �QAYLO vp2aHa1�]в�M1B�ׅ�pERVH�Af� �8l�-7�`�2��sE���RC\�ׅAScYM{aׅ�aWJ�'l�h�El�w1�If◁U�D�`Ha{5� gF�5aPZs5@
��6OR�`�M��Tw!��d���L001a��H9O���e �S1�,��OC�!��$OP���a.�F��䱩�`�2�PR�9aOU�sM3eV�RK5�U�X�1���e$PWR��IM�UIBR_�Sp4r�g `3�aUDlӳ3S�V	�eQ�df��$�H�e!f`ADDR
��H!GO2atama����R���g Hz�SE���壬e�ec��ep�SE?��bQyS����h $���P_Dq�����bP�RM_R��HT�TP_H�i (��OBJ��mb��[$��LE>3's>�j � |�b��AB_c�T#{rS�YP�s@�KRLiHITCOU�t���P ��P{r��l��P��PSSg�;�JQUERY_FLA�!�b�B_WEBSOC���HW���!��k�`�@INCP	Udr�O:��qH�Q���dR��dR�p�r�IwOLN��l 8z�yR����$SL���$INPUT_�!$�P��P�� ��}�SLA� m����مՄ�Cث��B�!IOpF_�AS�n��$L��Ow���1��"b�!`I������@HY��pX�1����UOP�o `�v���F�H�F�O����PP&c�P��@��O�ǒ���u�M�A�6�p lH CTA40BVpA��TI���E�&P ��0PS�BU IDC �r��?���P>�^q�:�?0qDЂ��+����N��| ���IRCAڰ��� r �my6ԀCY�`EA@�͡@��ҬF�&c�k�Rg0x�AA��ADAY_G�B�NTVAE�V�.�pȂk5:�.�SCA*@F.�CL��G����G���6�sr���l2����N_�PC⫠G��7�tЂ�Sޱ��Jr�G�>�p"�� 2�s ���6�up���Jr�LAB?1�3� 9�UNI�'�Q ITY���xe��R���vЂM�R�_URLT��$AL��EN�n�s�g ��Tv�T_Uk� s�J9�6�w X�����E��9�R����] �A�Ӂ��Jv���F�L9k���
Ӻ
��UJR��x ����FA�7��7<�D^{�$J7��O�B/$J8g�7P!�$p҂�78�c�8��f�oAPHI� Qq�z��D+J7J8�����L_KEd� o �Kt�LM��� y <��XR��G�ţWATCH�_VA��5@~�FvF/IELDhey����&��z R 51V>@¦K�CT��W�
�r���LG��{� �!��LG_SIZ�ut���� �����FD��I������� " ���S���� � �����" ��A�� ��_CM#3`���g�-F�An������T9(���2���@� ��������I��������" ����RS��\0  (�L)N[р|���p� @ڂ��,��s:YP�LC9DAU_E�Apt�|Tuk GH�}R�! �BOO�a�}� C7� `IaT�s�03�RE퐎�SCR��s8�D�I2�S0RGI"$D���+��T$�t �S[s�W� ��N+�JGMTMN3CH� �FN��W1K}��{UF��0n�FWD�HL�STP�V�Q �,� �RS�HP�(�C�4��B+�=P0T)Uq�/��>a�d@��Gm�0PO�'`���i�sOC��v�EX'�TUI{I��ĳɠ��4	1E@3yd��0G���	c����0�NO6AN1A ��QD�AI9�ttt��EDCS��c�3T�c�2O�8O�7S��2�8S�8IGN���G���zm��4DEOa5$LL�A��A�T��~F�u�T���$��l�B�ä���A\aF��P��M��p�� 1�E2�E3��Av��!�0 �m{Qk3�����?��=Q�u� ����FST���Rv Ys�R0P _$E$VC$[[�p3VFV ���� L4�F��P[�=�0#����Q$eENp$d�%6�_ � �p- p`�� �S ��MC-� ����CLDP����TRQLI]���	i�TFLGR�P�a+cr�1D:�+g%�LD+ed+eORG��/!>bU�?RESERVU��d��c�d�b�T�c� �� 	e/%d+eS�V 	`�	na�d>�fRCLMC�d�o �oyw��a� M�p���Ѕ��$DEBUGMASI��	äQ�uTu05�E��T~Q�MFRQ�Ŀ� � ��H_RS_RU���Q��A�T%FREQ̒�Q$%0��OV�ER-���o��FA�Pn�EFIN�%�Q��]q�T�q�d� \8���q��$U�@޲g?�`G�PS�@
��	�sC~ �c�W��sU��bq?( �	v�MISC.Ո� d6�ARQ��	f��TBN� ��&1ˈAX�R��·�EXCES�ºQ��)M���щ�����T��R��SC�@ � H۱_����pS�����PJPT��g� &�i�FI�����MI�� � ��Po�^H R�CT�Ns�ȖO"ҚAҚ��ԐC��u�^ԐUSEDw O�@TЏ�PX������@����^P)�/�+eR� ��pSZ��B_FR0�`T��\�Z_��^�CCO>� PHqK��a�A�h�cuB_���LICTB� QU�IRE=#MO��O���)�5�L�PM�Ŏ �P���r⛣�b���NDK���Џ�4+��9�Dx�GIsNA�DRSM\�S��0ё�S#��P�'�PSTL�ѐ �4��LO̐�DRI���EEX��ANG�k2k��ODA�uő��5�=���MF m����v�I�RA�U&Ŝ( avSUP�U4�F� �RIGG� � ��`�S'���S G&�T��Rn�P~ȀP��r��#mqPGW�T!I/��@��(�M\�Qr�� t�MD��I��)�ƕ0�q�H8ϰk��DIA���ANSW"�mA�!j�D})HqOR�b\�`�Д ��U��AVB��`k�j�_Lp�ѕ ��@�C��Np&+�����P�� 4����P��KEI"����-$B�p��zPN�D2r�a�2_{TX�TXTRA�341�%r���LOw ��1�$�G�T�F�.�|�g�_�ڲRR2>���� .W�[�A�a d$CA�LIĀ(�G�1��2΃@RIN���<$R��SW0t��%swABC��D_Jิ�k���_J3�
��1SP��r�k�P��-�3,���vPk�B\�J%sl��b�aO.A�IM%p��CSKP j��> qs��J~���Q����������İ_cAZ�bh���ELA<g�qOCMPҳ���J���RT�q)Y�11�i�G�Ȁ1�K40:Y
ZWSMG ��v3tJG�PSCL����SPH_�0����`k���RTEIR���S0��_�0
�Q�AS���sDI�23U��kDF^P�LW7VEL	aIN�R0&_BL�0k�.���l�J3LDMEcCHPB%r4�IN� �q���|҂�2�ҁ:sP_�� �����Ч?�����УDH�3഑�v@�$V��R��41$�v �q�r��$�a�Roӵ��H �$BEL �w�_ACCE4(�S'H%qa ʐ_� �q��iTJ��C*�EX�RL6��&c�w'��w'�.�W)�'m#�'36�RO
�_�A!"� 1�u�u�W!_MG�sDD!1��rFW�`��]#�=5m#X"28DE[;PoPABN�'RO� EE2�A�?	`��APOqO�X!^P�_��vbSP�pCTR�4�Y}03 �a yQYN���A���6����1Mwq�ѭr0O ��CINCa�̱Z2A4˂�:G��́ENC� L���k��!X"Ʉ+�IN��BI6��E���NT|ENT23_�r�CLO�r�@�pI�U��Fj��\�Ȑ@ia�C��FMOSI&1y���1�s��PERCH  k�q� .Wұ9S���B�3t��$�5)���A�"�UL�4��t����EpF��J�V�FTRK��AY[�(�O��Q�"�ecͰ/S�HB�pMOMc�˂O��`��T��Y3��c�#�2��D�U��7�S_BCKLSH_C�"�ewp V�p�3j��caB�jA>��CLALM�D}q8>`��eCHK����>�GLRTY���Ӑ�D��?���_�T_UMps=vCps/1��Us�pLMT)�_L  nt+�ywEs}�p �{rp�%�u�(>�aA��P�trXPC?QrXHpI�۠%5=uCMC7�\/037CN_��N6�L4�t�SFE!cYV�2���wG�	��"x��CATD~SHþ�34 iF?�xaxFX�7�X�L f"0PADt8B_PCu'c_�� f"P��c&�uJA�T�a��?�|'��TORQU�0 /� Sii0��R�i0��_WVe�TU"!��P#��#��I��I��I#F尜�s�����+0VCW 0�1Wd��1%�#09���+�JRaK%�j�]�u�DB� �M��u�MP�_DL!�RGRV����#��#��H_^㈣� �תCOS�1 �LNl��(�� 	�v @	�ۑE�3�����Z�V��MY������|����THET0�ENK23#β#�[CBӶCB#C��AS����۔�#��ӶSB#$�޵GT	S��1C0� �O�x_Z�B�$DUp@�W£�5��DQnQY_�sjANE���!AK$t;	��±AƵ�����֥��LPH��§E��S(�@�3� @�B���Q�j�T�q���EV�V� )�V8�UVE�VS�Va�Vo�V}�V��H�*�0�P(ݭ�G�E�HS�Ha�UHo�H}�H��OܥO�O��'�O8�O�E�OS�Oa�Oo�O
}�Oq�F���O�3��T��SPBALA�NCE_���LE6;�H_ƵSP�$���3���B�PFUL�C�������B��1=�=UTO_pu�T1T2	S"2N �a^"�@3�7a���(�"N#RaT�PO� `!>��INSEG^"�A�REVX�@�ADI�F�U�1���1��pOB��a��dg�2u��@q��LCHgWAR}2�2AB��feo�@��
AqXsX
aP�t)��� �� 
*��L!yEROB"PCR�"l��� �CJ!_�T �� x $W�EIGH@i@$�ӥ)�IA�@IF��1;0LAG�2�rS��2� �2BIL�O1D@`�@�STd �P��`��1 ���
���
]@J"�1��  2��D�DEKBU�L� "~�OMMY9�%� N���m$i@$D�!IQ�$W $���  _�DO_� A�� <�'& ���1���B��N�C�(_��@�0 "O�` _�� %\pT�@ĈA[qT�O$� TI�CK�� T1� %3�`(0N"P �#"PR�`�1�:5�F5� _PROMPCE�? $IRk��1pp�2�P�2MAI��h2A	B�5_��3� a@R��COD�,#FU�0�ID_�AP�5� {2��G_SwUFFې �4�1�152DO=7x >5�=6GR��D [3&D�1E�=Ev�DԞ$6 ��H� _F�I+!9�CORDf� �_"36�r��B�1� $ZDT��5� �%�4 =*�L_NA�!(0|�B:5DEF_I�H �B`6TF5�96$9602SF5@U`6IS��l� �!��94ySF3T�"]$4=��r"D �b��T,#Dh�O��"LOCKE��C:?L?0^7{QB@UME�B D2SD@UD�R&Bc %ES&DPT&B&{f{Q 1C� �1E�B1E2S1C�g�eH� P� iT� �uQ��� W�X�e�S?���TE�a�$ߣ �LO�MB_r/w0�V�IS��ITY�A�$�O�A_FRIWs� SIuQYq��!R%0�w00�w3E#��W\xWh{��^vn�_�y;AEAS�;B5��Vtŀ�P�2�v4~y5�~y6�ORMULwA_I���G�G_� h S.7e%COEFF_O1�o r�1C�G���S�~"CA���/�#!�GR�� � �G $�PF�"X� TM�W܄�U2�S���#ER� T�T�D6 7�  ��LL<D�P�S�_SV�TH��$v6 ���G�6 �{ ΂SETUuSMEA�0�0��!|�B�� � q�] g @����µ���Q���B(0�Q�Q�T���qFB�f1�PA�Q�P����� �0�REC�A���!S�K_��� P~�1_USER/��N�? s�N�/VE�L�N�? v�j��I��@� �MT�!CF}GD��  *0z� ONORE��� ���� ��� �4 ���X�YZ�C�@ J#	�ʠ_ERR�� ����!�0���2!�:���� BUFI�NDX��M�OR� H�CU��!_��1�A��<��A$Lt�AOQ�C�@ ��GĂ�� � $SI`;��p�0{R�VO��<���POBJE�����ADJU�"´ѰA�Y�AɳD��OU��@�_��1�B=�^�Ta .�v�-ǡ"DIR2�:�� ��ziGDYN�ry�v�T ���R^q� ����O�PWOR�� ��,� SYSBU���SOP��4�_���U�ˡ P�P���ŃPAQ������OP/@U����)"�f!�IMAG$���&�"IMw�@�I�N�p�?�RGOVCRDk���R��PЀ>�i� �`�S��L��PB�� ��PMC�_E�@4�[!N��M���f!_"1d"��k�S�L��E�� ��O�VSL�S�bDEX�QNP �2g ��_k��a@l��a@"�7�2�_"W�CZ�@�xf�4�l�_ZER��q�҃�D�� @נ4��3O�0RI±D
��0������*ܰLD��Z�T �ATUS��u!C_TV�C��B���������Se!���@E�� D�!���s�v3�0�A?�$���XE���\�p�;��㲠��cUPPoQPX�0�.��]$3��7���PG�����$S�UB��3]a����J?MPWAIT��'�LOW�1����CVF�1+0RXK���&CCi�Rm��2_IGNR_P�L��DBTB P�sQBW�0U��UL� TIG�j0IOTNLNS�R����R]pNj0��PEE�D��	�HADOW ��ʰE�����PSPDD�� L�A'�P"�0CUN���.��Rw��q�LY�@�  ���P��D���$0���f0� LE��� �PA�P�����I�P�~�S�ARS�IZ�4�@�CMQܰO8>@�9�ATT���8-����MEM�"f!��TUX��}�L��0��� $���aS�WITCH	�!W�ͰAS���A0#L�LB~�� �$BA+�D�S�BCAM��[Å)��w #J5����"6�&Y!_KNOW��"k��U�ADz(��-D�Q��)PAYLOA���`3_D�7��7�Z3L]aA��>PL�CL_� !@}�D2�!��Q4��_6Fi9C�?:��B4[��I?8R�?70�[4Bd�p�Jq��1_JI1:i���AND/�
�`�4I2]19��qPLh ?AL_ �= -P���!��<pC�D3�E��J3�0F�{ TU�PDCK���rR�CO��_AL3PH CfCBE��(�� O2L������ �� �� ?D_�1:224D��AR�c��H�E�F�C��TI�A4Y5Y6�MOMq�S:S'S:S4S��B% ADS^V'S\^V4SPUB��R?T �U'S�U4Rq�@G@���  �M,2� v1!A���� e$PI m���CZ�7i`�'9*iIkIkI+c�T �\f��\f����\Bpg�Wª��HIGL# �&�f&\ K���f�c�h\�i\&SAMPk�d�t�gs8&� �3 �Fq ��z�Ut��_v�@ ny�@z�����P]u�q�b]uIN�|�p�c�x �{�t&�z�x�t�{�/GAMM�uS
���$GETW�@���iD�D��
��IB����I�$HI�_�[�D�z���E����A������LW��̆Ì��������B�f� AC��CHKyг�ڐUNI_�`����B�H �q�uY�RS��|VX�GC� �$BH �1���I��RCH�_DX�����G��L�Ev�Z���嘩H���>� MSWFLV�Q7SCR��10���	SN�Wr3��:�|w��PnyN�]�PI3}A�VMETHO}�X�����AX��h�qX� ���ERI��Jt3C�RB�5	�a"�@F4�q\s��ks���LĐq�O�OP\q��0�kq��APP��F�И4��U�@��sRTբ�O �0���a����T`1���T`஺+`���)�MG��,&SV~�PD�G� ����GRO� ��S_SaA�!��ū�NO�@C���D�b��O? %?1h�o�W`�"_e���CDOA_�� Uv P��u�h��g��hט���H3 9�0 M��U� � ^�YQLc�1�w��S�2Q��b�(����1���nӽ1_đC�Z�M_WA��� �w����Mj ��d0��A3A)�	(����PM�~�R� � $Y�Dm��W"�n�԰L! 51"��D �D �D �4D{ ��N� d�C#��J�pXjO�C�qZ���P0 �T� ���M��W�T�f�xϊϜ�PP��ّsL�A_��� |SA���:Yl� 'Sl�4S�Z����-Z�R!\�*%P���t�60P�P��PMO�N_QUp �{ 8�QCOU��n�`QTH� HO[�n HYS�ES�"F UE µO5$�  ? P �|�3��RUN_TO��q�D �b�P� P� �`C��/���IND}E��ROGRA���' o�2��NE_NO�`IT�Q� D �INFO��� �?!�
�m���OI��� (p�SLE�Q�f��e� ���OyS2��� 4��ENABN�^ PT�ION���ERV�Edb[ra��3GC]F<� @ J�Ь�qh�h�R��\n�R�PEDITN��� �/��K�Qj�c��E��NU���AUT.��CO�PY�Q�`,ra:�M⊁N +*�PRU�T�R "N�OUC�a$Gep$���RGADJ��� -hS@X_��I͓��(�&���&W�(P�(�М&�c� �N�0_CkYCN��#NS89�P��`LGO7�s@�NYQ_FREQ�RW�p�f-1SIZK8�LA��$1�!5S�p�eCREo���8��IFa�NA q�%k4_G��STA�TUS�VMAI�LrbA�1�LA�ST�1aA�$ELE�M<� �9�FFEASII�KrD� t��2���F٢�pn�I� l�$2�a���&KBAB2�@E� �`9V�1cFBAS�BdE�n��QU�`�`'�Y${A�GRM�PREC �qؐ�C���`��1�D� �5�S�[�	~"B 2� �s ���tV�BW�B�Њp��ѡB3W�WߔDOU��ӔO��$Pݡ�@ОGRID�2B7ARS�gTYJ/r�pO����� QE_�4!� �RnTO��>9� � �����POR��S���SS�RV�0)�T�VDI0�T_e``#dr`-gT`-g4+i5+i6+i%7+i8a�F?�<��O $VALU�~C�DG�a9��� !E;��S�1�۠ANõb�1�y�12ATOTAL�_�4I@rPW3I|vQ(tREGEN&z;r��X�Hu����f���TR�C�2&q_S��w;pأV�!��rsdBE�3ݠB`���cV_H�PDA8��p�pS_Y6����>6S�AR��2�� h"IG_SE��p�R�5_d �tC_�V$CMJ�C�T�KDEE��b�I:��ZS�-�N1�FB�H�ANC� p��AG�2A3�qIN�T`�!��FZ��M�ASKʣ�@OVR ����ݠ��1��WV�AߠzT�A�_'Fd{>�V�PSLG%��a� \ �?57���p�0S���4f�Us�V|��s��7a�UP�TE���@�' (cq��J3�.N3IL_MM4�VQB۠��TQ�𖣷R�@C����V�C-��P_�'�7�MN�V�1M�V1[�2j�2�[�3j�3[�4j�4 [�����ޣ�ޣ����;IN��VIB�'������2�2#�3*�3#�4�4#��� 6�O�2���D`�Q`�����PL�0TOR ��INƵ��R���L��T $�MC_F  5�B��L ����pM?�1I���OS ]���f���KEEP_H/NADD �!B�h@L�C�ᐐbĮQ�t�c�O��A� ���p�cë�c�REMz�@bĺ1�R�Ŷ���U�4�eb�HPWD  ;B�SBMӁ�P?COLLAB���`he�qq2� IT0��&"NO�FCAqLE����� ,���FLK��A$SY�N��`�M��C@��~�pUP_DLY��=�ODELA�л1Z�2Y��AD�����QSKIP$�� 	��Pb Op਒(���P_b ��ד ���  �׵ �s �D`��Q` ��^`��k`��x`�څ`z��9�!�J2R� *���AX�@T'3�� �A�� >¡�>�μ�RDC�aT�� %��R�˸R`1ɺ8Ȳ
TRGE�4CгXRFLG���ŐsSWX
TSPC���!UM_��ؓ2T�H2NRQk�� �1� ��ED|�Q8 � D� x��:�l@2_PC�#��S���A.0L10�_CL2䱅�́ �� b�'`����F(�@������ ��+U���г+� �b9�lC���������~D�ESIG��'UVL�1��1��Hs10��_DS�(�G��pv  11�� l3�`i���o�F&�AT��@q$]Q07�'+$��  ������HOMME ��2�������! �3��DVh�z�� �4������	//S U�5��>/@P/b/t/�/�/36���/�/�/�/?? )��!7��8?J?�\?n?�?�?�'8�逵?�?�?�?�?O�S|���  �A��Pp6�3��E�T�� T���D	v�CIIOՑ�IIp@5�OB�_OP�ESr�C��POWE��� ��@_п�."t ��Z�BR$DSB�f�GNAOs��Chq�a�!M���Z�|CIk T_SPE%�-z�MD�W_�Q�dy��DBG_\@PU�����SEq�̀� 2�4C=�3Sw232�E� ����7Eo���ICEU�Ss�U�ARIT��qqOPB.ЭbF7LOW�TR�@r���P�aCUV` �a�UXTҁ�a��ER�FAC;d��U�`��2SCH��� �t3����QH�@�$L�p�pOM���A�8  t��UPD���f�qPT�@Y�EX��4x�c!�FA�e����qfq � h�цp�� (�AL� �3u���:R;�  2� �S��~�@�	� �$X�z��_�GROUQ�sT\ ��vDSP��vJOGLI�cF����,a7�N������ސ�fK�`_MIR��q�T�MT��A�P��c�*�Z�`�S�Yq�t�]��@�BR�KH�avl�AXI~A  f�@�q��r�ρТu�BSOC��v��N��DUMM�Y16,�$SV��DEQnSFSP_D_OVR.���2�D؂�sOR�P@�N���Fv���pO�V�uSF�RUN����F8��a�sUF�RAN�TOldLC1H�Ҥ��OVׄ8��pW- ��sy�P���r��_8�ϰ @E�TINVE$PKAO�FSǐCSp��WD� ��������R#�ÀTeRO�R(�FD�Þ(�MB_C4��B� BL~���q0�6��qPV�adB�` ��2�G1�D�AMB�$�0�`r�����_MH��b<��C��T$����q>~CT$HBK�a/�ءIO_E�Q��PPA۪�����x��R��DVC_�P dCI�q`RI�҆a`�1h���`�3h���"���`�pׁUdC�p�FCAB��^B[�"��h&�k�h�O�UX/�?SUBCPU_R�pS�����Z��`���I�Z�?R��$HW_C� t`���N��qN@pNp�$U-��z�t�m�ATTRqIEЁ��pCYC���ұCA���FLT?R_2_FIqCsY賳fV��P�{CHK�_�`SCT�F_�m�F_w� ҉�FS8eQR�r�CHA����pA�Q�{b@�RSD��`bQ��s`QP_To�0? ���q`EM�@��EMn�T.��Np.Ҽ�Ӷ�DIAGuR�AILACV���M�pLO��f�<�'$PS�r`B ������PRJ�SZ�& ��C<�C 	��FUuN��aRIN��Z�Y@��?�pa��S_�pu àh�@Ѥh��-�ѤCBLCUR�}��A������D�Ax�i�����LD@�`ˀ����qr� ���TI��}�Np$CE_RIA��oRAF�P�SG�[ L�T2��Cs��C��OI��DF_L��@P��as`LM�SF>;HRDYO�ѐRG �Hb��Y@��>��MULSE�����Ǽ�s�$J�J�����FAN_AsLMMWRN!HARD`@�ffs�!2Vaz�R�_��/��AUR�R3ԇbTO_SBRU��p�
�m�>�G�MPIN�F��������REG`FNV�`�Sb�5DPN�FL_Ž�$M�����c��Np(/C�P� ��FdA��PӐa��@;$qA$Y�R�a�}r�S�� �7�EG&P�sˀb�A�P�D��25������D�AXE�wR�OB�zRED�vW�R�Pk�_���SY�h��Ϡ&S!'WR1I�P�M�STOP�s(�`l��Eo��@�6��f�pBa ��h&�7�ӝ�OTO��@Y�ARY�s�"�ј���B�pFIM��s�$LINK��GT5H�"
pT_^#����8���!XYZt�b�*9�&OFFŐP�"�P� �(� B�p�4�D4��m`�`E3F�I��^7K�nSÄ4��t_J,aNr���#��[ w$�*30��9`�ȕ1���2C#Q4�DU��³�3%���TURB X"�E�!�X0 `�7FL� l�̳��$@5d)35�Ғ W1��@K�pM/���6�������cORQ�ֺqn�8��J�O N��E���q�N�DOVE�A�RM�` �Aj
Up
Uv	Va`WαWpTANE� �!
QL�Q�A�IP�� QU�AW�Up�U.S��qER�qr�	 �E���Dp��TAQNp�a5`�ҫ'��׶��AX��Nr�ᝰV��"+e ��7i��7i��6j�6j q 6j� 6j� 6j06j1�06f��3i��Ci�� Si��ci��si���i����i��i��i�a�iD7EBUE�$@�L0��tqڒ�"AB��ء� ��CV͠D� 
 �rq�r�u5��w���w ���w��wq!�w�!�w �!�w1R��0L��"E3LAB[2�EA�N�GGRO���2E��B_�ѸVM$��U0� �l����E��y��ANDr@ ��T���%�Qy� ��M^ ��������� NT, ��+�VEL��eT5���=����E3NAc�� ��$��ASS  O�������3 x�ʐSI����w��㆔��I��������AAV�M, K 2 ��� 0  �5�������%� %�	 H�9�\�����J���n���8�����G���0���АBSQ�� 1��� <�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e��nL�MAX�� h��5�  dz�I�N����y�PRE_EXE������D����АIOCNYV*B�� ȑ�P��p�0��1��IO_��w 1ݛP $͠��r�]��Z��?� h���}����� ��1CUg y������� 	//-/?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ����	��-�?�Q�c�z�L�ARMRECOV� �����6L�MDG F�Q k�LM_IF F��h��"�4� F�T���wωϛϭϾ�?, 
 ���πb�n��1�C�T�$ ��x�_ߜ�[�����������s�NGTOL�  �� 	 �A   >�P�z�P�PINFO Ż Ķ�������  �»��者 �����6� �2�l�V� ��z����������� (:L^p������غPPL�ICATION �?-�����ArcT�ool  
�V9.10P/3�0O��
883340-F0S@�105-"4�7DF1(�N�one�FR=A� 6p�_ACTIVEp�s  �7�  ��UTOMOD ���5��CHGAP�ONL$/ 8#O�UPLED 1�� u y/�/�/��CUREQ 1]	�  T�)�,�,	�/	5� 4����"_AR�C Wel���AW���"AWTwOPKS6HKY? ���/�/�/?v?�?�? �?�?�?�? OOO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ����(�:� L�^�p���ܟ����ʟ �� ��$�6�H�Z� l�~�د����Ư�� ��� �2�D�V�h�z� Կ����¿����
� �.�@�R�d�v��Ϛ���Ͼ������̹%TO�(�/#DO_CL�EANE/�|�NMw  -� �/������� ��.DS�PDRYR��V%H	I" ��@��~��� ����������� �2�8D�V��MAX� c��1T't�Xc�sp"|s�PLUGGc �d�p#%PRC5�B�����m�_���Ox��>��SEGF<  ^0.7�߶�~������1LAP [�n03 2DV hz������>�TOTAL����_USENU[ h+� I�M/2� RGD�ISPMMC^0z21C+3�@@�"�h$OY�{�I�RG�_STRING �1
4+
��M- S�
�!_�ITEM1�&  n��/??%?7?I? [?m??�?�?�?�?�?��?�?O!O3OEO�I/O SIGN�AL�%Try�out mode��%Inp�@Simulated�!�Out�LO�VERRX� = �100�"In �cycl�E�!P�rog Abor��C�!�Dstat�us�D�@cess� Fault\A�lerT	Hea�rtbeaSgCH�and BrokeZEWOY_k_}_�_�_0�_�_�_�__��+ _��/�_9oKo]ooo�o �o�o�o�o�o�o�o�#5GYk}�_WOR: �+�q)o�� ���%�7�I�[�m� �������Ǐُ���8�!�3�PO�+1Q Y��{B�|�������ğ ֟�����0�B�T� f�x���������үT�DEV\���p��$� 6�H�Z�l�~������� ƿؿ���� �2�D��V�h�z�PALT m���{��������� �#�5�G�Y�k�}ߏ� �߳�����������GRIy��+E��� m����������� ���!�3�E�W�i�{� ������3�+ Rm�� ]���#5GYk }��������1CU��PREG�Ύg�� ���/!/3/E/W/ i/{/�/�/�/�/�/�/��/[M�$ARG_��pD ?	����<1� � 	$[F	+[P8]P7�[Gq9�/0SBN_CONGFIGj@<;�A�B��1�1CII_S?AVE  [D�1��3/0TCELLSETUP <:�%  OME_I�O[M[L%MOV�_H�0	OOREP���ZO%:UTOBA�CK�1<9�2�FRA:\{ �eO{�0'`�@�{�H� �K�0� 23/0�8/13 15:_18:50{r8�{_-_Z_Q_�L�� z_�_�_�_�_�_�_{��_)o;oMo_oqo�o o�o�o�o�o�o �o7I[m� ������!���ׁ  �A_}C_\�ATBCKCTL.TMH�`�r�����\��oKINI���E��5�1z@MESSA�G�0ρ�1D0ڋODGE_D�0�6�5��O���wCPAUS�m� !�<; , 	�r0<5q��,		i����� ǟ��ß���!��-� W�A�{�e�����D�N�?TSK  T��O<��z@UPDT�͇�d��XWZD�_ENB̈́�:'�SCTA̅<1�.1WJ@�ODP�2<;�4W�)13-AUG-2P7:33P42O�� ˿ݿ奫3{��R���&�4�]�{7u�C�� . �� �9�fϚ���j�R�OBGRPҨ�AS�"�WEWE�Lp���k��6~��3:24:4���E	LAB��_2��{���9k�f���q�oߢ߯���5 �C 5 ��  f�����oAXIS�0UN���Ԧ�1��� 	 ��	 �� M����{(<;�V����B�C�1T��H�{��{V���K� �� - ����� �,����������0�3�MET��2�D鄰 PU�A��m@���@w��^@(��@�ߴAQj�?�%�>�E�=��i?I�>���0?�@��5�S�CRDCFG 1�<5�A ��5�2���);M�O{Q�9��� �����^� ?Qcu�� :'7}AGR=��2���C�NA#@;;	�}D�_EDˀ1���� 
 �%=-I�EDT-���m/����@!~BI/�څr2p_FB/�/  ���%2�/6K�/ F?7��+??�/�/n?�/�#3�?'?OK?]>��?KO�?�?:O�?�#4 �O�?�OO]>�O_^OpO_�O�#5O_�O�_ �O]>x_�_*_<_�_`_�#6o�_ho�_]>Do@�o�_o�o,o�#7�o Wo4{o]>{�o�oj�o�#8�[/ ��^=�G���6���#9��̏�h� �)���Z�l�����!CR�/"����X}r��ݟ$�6�̟Z��% N�O_DEL��GE_UNUSE���IGALLOW� 1��   �(*SYST�EM*��	$SE�RV_���ٗ�POoSREG��$£�ܗ�NUMŪ�ح�PMUC���L�AYO���P�MPALS��CY'C10$�7�!�%�]�ULSU�٭9�� ��Ls���BO�XORIɥCUR�_��حPMCNmV���10M�~��T4DLIB�����	*PROGR�A��PG_M1I%�O�a�AL/�n��X�a�B�ϗ�$�FLUI_RES�U=���ϯ����MR��������Wr?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ��������������%�7�I�[�6�LA�L_OUT ����#�WD_AB�OR>�g���ITR_RTN  �������NONST�O �� O�CE?_RIA_Id����0 � FCFG *0���9_PA��GP �1CU �����C;��i� ��C� C � Y(� M�C8� @� YH�  CX� `� Uh� p� x��� U�� �� �� �R�dv���?�H=E�ONFI���n�G_P߰1C 1�����/� /2/D/V/h/�KP7AUS��1��0 M�j/�/���/�/ �/�/?�/6?H?.?l? R?|?�?�?�?�?�?�?�r,M��NFO 1���S  �� 	�OO;�=@B�7��yO  ��'��Dd��8C��6����X hB�@��d��ðXD�̿73��¿W���3�gO�=C�Ǹ�CO�LLECT_=b+F��R�GEN/�p���R�ANDE�C��GR��1�234567890[W:ұ�SY_kV��#
 %}�;�)�_�_ ���_�_o���_�_To o1oCo�ogoyo�o�o �o�o�o,�o	t ?Qc���������L��5V��2��K ]9RI�O !DYQ�����Ώ������TR�r 2"�� ��
-���#��<��^Y_MORz�$w ��ŕ<Ařݟ˟���%����m{�%J��,�?���x�B;�K��;ѷ� R=�&�O������C4 � A����;�=}A{�Cz  B��$B�"  @�Ң��;�:dڬ���ARI=S'��?D�z�(���/�d���T_DEFz� �X�%J�������NU�S<��0��KEY?_TBL  �0�6B�	
��� !"#$%&�'()*+,-.�/dW:;<=>?�@ABCe�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������h���͓���������������������������������耇�������������������s��}!b�LCK��8	b���STA�����_AUTO_DOr��&�INDT���_T10�"�T�2o�V� TR�Ld�LETE�����_SCREEN� �kc�scU MME�NU 1)�� <o�|�D�UE#�M�� i�k���������� ��6���l�C�U��� y����������� �� 	V-?e�u� ���
��R );�_q��� �/��<//%/r/ I/[/�/�/�/�/�/�/ �/&?�/?5?n?E?W? �?{?�?�?�?�?�?"O �?OXO/OAO�OeOwO �O�O�O�O_�O�OB_�_�_MANUAL���DBc�j������DBG_ERR�Lj�*�D� �Q_�_�_n�QN_UMLIM��[����
�QPXWOR/K 1+��__o�qo�o�o�oS�DBT;B_�� ,�]ģ�4���o�DB_�AWAY�SD�GwCP ��=��1b�b_AL`��b�R�Y���ը��X_�P +1-��h�
No����|��f_ML�I�S�
{@{��sON�TIM�����ɼ�vGy
��\sMO�TNEND��[tR�ECORD 13�� ����G�O���u���
r��ŏ ׏鏀�����<��� `�r����1���)�ޟ M���&�8�ӟ\�˟ �����ȯگI��� m�"���F�X�j�|�� ���Ŀ3������ ��Bϱ�M�տ�ϜϮ� ��/���S���w�,�>� P�b��φ�q�߼�+� �����s�(���^� �߂���=����K�  �o�$�6�H�����~� ��������������  ��D��hz����bTOLERE�NCtB�QrpL��͈PCSS_C�NSTCY 24J?i��P�Or�	 );Q_q�� �����//)/�7/I/[/�DEVI�CE 25� �f�/�/�/�/�/?�?,?>?P?b?��HNDGD 6���`Czu:O��LS 27�-t?�?�?�OO,O>OPOv?�PARAM 8hy�8rwUbD�5�5SLA�VE 9�=�7_?CFG :�ObCdMC:\� �L%04d.CS�VaO"�c	_!�>AM 6SCH>P�1�PbNI_~_�G�bFnR��Q�_�Y�Q�@JP���S�^"��a�>_�CRC_OUT �;�-�afO_NOWCOD�@<hw�M?SGN =^�G��#M�16�-AUG-23 12:399P�Av`�3zf5:1�a�&? Wzz�i�a�bN�`ra�M��?Þ�j��a�n��CVERSION� ejV4�.2.11�{EF�LOGIC 1>^� 	�X�@�Iy�QY}+rPROG�_ENB<��6ysU�LS�w �6+r_�ACCLIM�v���C��sWRSTJNT�F��A�+qMO�|�QPb�tI?NIT ?�
^�v�A �vOPT�@� ?	6��
 ?	R575bCc��74h�6i�7i�50��t��2i��X��|%wF�TO  R���o�&vV�DEX��wd�riP$�PA�TH AejA�\�q����HCP�_CLNTID y?	v�C �[�Zß�IAG_G�RP 2D�I �> 	 �@K�@G��?���?l��>� �ٚ���8�ٜ5��� a�O�?ϧb�?> ��i��^?�Vm?S���ٙf403� 6789012�345����� ��s��@n���@i�#@d��/@_�w@Z~��@U/@O��@I��@D(��ٚѠiQ@�6TpX6P�� A�� � 9PB4ٜ� ٔR��iQ
Т1��-�@)hs@$���@ bN@���@ڠ��@?�D@+2�	���-�2�A�2�P�R���@N@I��@D�@>�y@9��@4���.v�@(��@"�\��������п�V�L�@Gl��@BJ@<z��@6ڠ0�`@*��$���@��&�8�J�\�V��=q@���F@|�@3�3@�R@-�?���?��`?�+�ϲ���������̑҂��-�@&�@�����!?�?� �,�>�P�b� t�V� �(�:��^�p� ��D��������x� ����6�H�&�l�~�� ��:���q�����Ѥ��x������Y�?��?�z���(�o5AF4� ��L4R� �(�@�p�8�Q��@-: I �m@����%�Ah.�=H��9=Ƨ�=�^�5=�v ��>��(�=�,v��,�^ �iQ�C)�<(�U�Rc 4�����ٙA@hR?0���"�� 0Vh4��t�8�����
/��>���y,"�R=�?��=��z<!(�o��G�T/G�(�@8U8U����(�$@9P���*��uB��J���B�B�?�B%�(��T$�/�.'�p5.�*11n,�\��=�-���c+�a Bk B��BC�A��@�Z?؟�?�iQ<�P  3�>��?y?�O��3P1����3\�N2�J�d��0�18��BDd�8C�3Q�>�V�?O�?6O�+�TOZBٙ�96���.�B�R�)O�O��O�O�O�O�O__�>�{Dٙ>�� ���'_u_��CT_CONFI�G EDo�c�eg�U�STB_F_TTS�w
�y��S p�s��V5`M�AU�p��rMSW�_CF�PF��  �)��jOCVIEWf�PG'm3���ן yo�o�o�o�o�oPrgo �o 2DV�oz �����c�
� �.�@�R�d������ ����Џ�q���*� <�N�`�������� ̟ޟ���&�8�J� \�n���������ȯگ,�|\RC cH`��R!����$�Y�H�}�l�𡿐�ſdSBL_�FAULT I��<h߱GPMSK��W�PTDIAG� J�Y�!�S���QUD1:� 6789012345O¬RC��W��Pb_�ϝϯ������� ��	��-�?�Q�c�u߀�ߙ߫�j�?���
�z��߂VTRECP(�:�
H�:�a���y� v����������� ��*�<�N�`�r��������������=gUM�P_OPTION�P���TR b�S﹝PME�UY�_TEMP  _È�3BQ0m 9�L1WUNI`�U�m�YN_BRK� KRo=fEDI�TOR��F�_~�ENT 1L��  ,&M�AIN LD_2�����&	LABW�E@&
*_-1A��T2���ֲ���� /�/C/*/g/N/�/ �/�/�/�/�/�/�/? ???&?8?u?\?�?�? �?�?�?�?�?O)OO�MO4I� MGDI_�STA�+am�N�CsC1M'k �P���O�O��
��d�� _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o&�o �o�o�o�iQ�o" 4FXj|��� ������0�B� T�f�x��j�o����͏ ߏ�o��'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uϏ�}ϫϽ� �������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� �ϙϣ����}����� �!�3�E�W�i�{��� ������������ /ASe��� �����+= Oas����� ��//'/9/K/]/ o/��/�/�/�/��/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgO�/�O�O �O�O�/�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oyOko�o�o�o�O�O �o%7I[m ������� �!�3�E�W�qo�o�� ����Ï�o����� /�A�S�e�w������� ��џ�����+�=� O�ɏ{���������Տ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�s�}� �ϡϳ�ͯ������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�k�Y������ ��������)�;�M� _�q������������� ��%7Ic�u� ��Y����� !3EWi{� ������// //A/[mw/�/�/�/ ��/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKOe/ oO�O�O�O�/�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCo]Ogoyo�o�o �O�o�o�o�o	- ?Qcu���� �����)�;�Uo G�q������o�oˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�M�_�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+ϥ� W�a�sυϗϱ����� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�O�Y�k�}� ��ϳ���������� �1�C�U�g�y����� ����������	- G�5cu���� ���);M _q������ �//%/?Q[/m/ /5/��/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO 7/I/SOeOwO�O�/�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'oAOKo]o oo�o�O�o�o�o�o�o �o#5GYk} �������� �9oC�U�g�y��o�� ����ӏ���	��-� ?�Q�c�u��������� ϟ����1�#�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ��� �)�;�E�W�i�{ϕ� �ϱ����������� /�A�S�e�w߉ߛ߭� ����������3�=� O�a�s�ϗ����� ������'�9�K�]� o��������������� ��+�5GYk�� ������� 1CUgy�� �����	/#/ ?/Q/c/}s/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�?��?O/ �$EN�ETMODE 1�N~%� W + + &%�HOZK*@RROR_PROG %7J�%%&�O�IxETAB_LE  7K�/��O�O_WxBSEV�_NUM FB  �AA=PxA�_AUTO_EN�B  dE?CuD_;NORQ O7KYA}<R  *��P���P��P��PHP+��P�_�_�_nTFLT9RZ_lVHIS9S)!�?@g[_ALM 1]P7K �&$�\% +�_no�o�o�oȶo�o�__2RtP  �7K�QZBz*@T�CP_VER �!7J!�O�o$EX�TLOG_REQ�f�eY_sSIZ\hZtSTK�y�U��\rTOL  �)!Dzb�A= Zt_BWD�`�p��V�q_B�sDI�q ;Q~%�sXD<)!�{STEP��|*@0�OP_DO��(AFDR_GRP� 1R7I�Qd 	���Z@��n&����c?���$,MT�� ��$ ����ن�������Bؘ��CF��B���rCP�B�ϘB��H`�A��0�A��B��]�B)�jA�?WA������ r�]���������ޟɟ�  @�?�A���>(��A��`�
 K_�A�	�)!A��g�Eb؟ҟw�b����*�@7���@�33K@�Ǡˣ�@¡�毄�����F@ 5�E��@�5�%���L�FZ!D��`�D�� BT��@�����?�  ��#�6������5�?Zf5�ES������E�K$FE�ATURE S�~%�p^AArcTool ��)"Engli�sh Dicti�onary*�4D� Standar�d#�Analog� I/O"�A5�e� Shiftw�r�c EQ Pro�gram Sel�ect��Soft�par�ǝ�Wel�d��cedureys���Core����Rampingn_�uto��waпUpdate(�m�atic Bac�kup(�V�gro�und Edit� �-�Camerazr�Fv�Cellr��{�nrRndIm�[Ӓ�ommon �calib UI�����sh������c��	���ne�	�t%y��s����nt���Monitor=��ntr�eliayb��)�DHCP����ata Acq�uish��iag�nosR�o���oc�ument Vigewet��ua���heck Saf�ety��-�han��� Rob��rvB��q!���)�F�s���F���-�xt w�eavS�ch%�x�t. DIO��nsfi"�|�end.�Errs�L���i�%s��rm��� �p'��FCTN Men�u�����TP I�n��fac�-�G�en��l��Eq 9L��8igE'9�m�p Mask �Exc*�gr�HT|% ��xy Sv����igh-Spe.�Ski�ԍ�����mmunicQ�o=n��Hour ��x��s�(connX��2�ncr' st#ru>��
!e����J��-�KAREL Cmd. L� �ua�XRun-;Tiq�EnvN���:�+U�sS�S/W�*�License������Book(System)'�MACROs,��/OffseZ�M�MRm�i���Mec_hStop��t��D���i���1&x.��o�S�D.od��wi!t��g(i���.�ƅ+�Optm�/#��f�il��'g��ulti-T  �+��ORNTBASE� Fun+-�PCgM f"8(�Po��x� �I=Regi�r��,6ri��!9~9�p�Nu����8��Adju� �>���=tatu}1�?��,ŷRDM0�ot;�s�coveD�)Eea�� q�Freq Awnly��Rem' ��nR�)E5B5�9�'ues�ńGo��r ~)�SNPX b�v#�SN% Cli���N��P rC��OU� �8$P�Eo�t ssag յE���Ob!p 0��V^/I&>]UMILIB�_`R?P Firm9�p^�PAccn�v�T�PTX��^Teln���_aQ��q]or��@ Simula(r��!fu��P8�XZ�mЍ�#&��ev.�]U1�ri��_U�SB po����i�P��a��fR E�VNT�o�`nexcept.�j@W4�e,j�P�VC��r��-(V��.r�_?u�K9{�S�@SC�UqSGYE�|uUI&�W��<8�|b PlF�~ 5���� (���������6�uZDT Appl�'��f�s��Grid9Apla�ym�mPZԇ�R%r.�R�����F� A�2�00i��c�lar�m Cause/�h@edE�Asci=i��Load��1�gUplG���yc��`~�0�`� RAe`x���yQ�NRTL�_�4nline Hel��-6',6{0x1���tr"�64MB� DRAM���FCRO �����c� PB:� .'�mai���K��RR�6L��Su�p�b�!}9à��} c�roL4C�E��9vrt�4C&���z�.� @�m�d�v�������ٿ п����3�*�<�i� `�rϟϖϨ������� ���/�&�8�e�\�n� �ߒߤ����������� +�"�4�a�X�j��� ������������'�� 0�]�T�f��������� ��������#,Y Pb������ ��(UL^ �������� //$/Q/H/Z/�/~/ �/�/�/�/�/�/??  ?M?D?V?�?z?�?�? �?�?�?�?O
OOIO @OROOvO�O�O�O�O �O�O___E_<_N_ {_r_�_�_�_�_�_�_ oooAo8oJowono �o�o�o�o�o�o�o =4Fsj|� �������9� 0�B�o�f�x������� ȏҏ�����5�,�>� k�b�t�������ğΟ ����1�(�:�g�^� p���������ʯ���  �-�$�6�c�Z�l��� ������ƿ����)�  �2�_�V�hϕόϞ� ����������%��.� [�R�dߑ߈ߚߴ߾� ������!��*�W�N� `���������� ����&�S�J�\��� �������������� "OFX�|� ����� KBT�x��� ���///G/>/ P/}/t/�/�/�/�/�/ �/???C?:?L?y? p?�?�?�?�?�?�?	O  OO?O6OHOuOlO~O �O�O�O�O�O_�O_ ;_2_D_q_h_z_�_�_ �_�_�_o�_
o7o.o @omodovo�o�o�o�o �o�o�o3*<i `r������ ��/�&�8�e�\�n� ��������ȏ����� +�"�4�a�X�j����� ����ğ����'�� 0�]�T�f��������� ������#��,�Y� P�b�|���������� ����(�U�L�^� xςϯϦϸ������� ��$�Q�H�Z�t�~� �ߢߴ���������  �M�D�V�p�z��� ���������
��I� @�R�l�v��������� ����E<N hr������ A8Jdn ������/� /=/4/F/`/j/�/�/ �/�/�/�/?�/?9? 0?B?\?f?�?�?�?�?��?�?�?�1  ?H541�3A�2FR782 G5�0 EJ614DG7�6 EAWSP,G1�[GRCRPH8\FT=UgFJ545DH[F�VCAM ECLI�O�FRI�GUIFz,F6�GCMSC�H^gFSTYLDG2�FoCNRE,F52[FwR63+GSCH E�DOCVLVCSU� EORSFR86�9DG0OG88FE�IO�FR547FR{69[FESET�G:rGJqIWMG�G�W�MASK EPRX5YX7 FOC�F�P�3�H7F�PCH3fJ�6BH53{VHEhL�CH�VOPL�VJ�50/fPS�gMC�fG�`�W55OFMD�SW�g"gOP"gM�PR�F<PSh0CFO�RBS fCM�G0�w�POG50Sg51֣G51Ox0�FPR�S�W69fFRD޻FFREQ,FMC�NVmXH93CFS�NBA�GFgSHL�BVM�w<P3WNN�_h2CFHTCgFT�MIV4@{VTPA��FTPTX(�EL��v�`{W86G4@FJ�95�FTUT#g9�5fUEV�VUE�C�VUFR�FVCuCψOFVIPVwCSCW�CSG'VraPI�hOFWEBgF�HTTgG62WWI�O�Ry�CG:�I�G�IPGvIR�CVDG"gH75��FR66��7�WR*Mz2/fR]j4f���OF�@FNVD�VDu0��F�ALO�V�CTO�GNNfMv}xOLXEND,FLڇFVR�E�8�� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿���  H5�41��2#�R7�82$�50$�J6�14T�76$�AW�SP4�1s�RCR�d�8t�TU��J5�45T�s�VCAM�$�CLIO��RI���UIF4�6��C�MSC4܃�STY�LT�2��CNREv4�52s�R633��SCH$�DOCV��CSU$�ORS^��R869T�0c˻88#�EIOC�R�54C�R69s�E�SET�˒�J��W�MG$��MASK^$�PRXYd�7$�OC�`�3��C�`��S�3��J6R�53���H�LCH��O�PL��J50��P�Sb�MC��p�c�5=5c�MDSW����;OP��MPRڠ�z�0S�ORBS��CM#�0`�c�5m0�51��51c�0��PRSS�69���FRD��FRE�Q4�MCNT���H{93S�SNBA$�^�SHLBT�M2��Г�NN#�2S�H;TC��TMIc�@����TPAC�TPT�X�EL�
p���8�B�@�#�J95��T�UT��95��UE�VS�UEC��UF]R��VCCc,O��wVIPc�CSC�'CSG����Id�c�wWEB��HTT��]6��WIO�*R��CG�+IG�+IP�G#
IRCc�DG���H75��R66��;7B�Ra2��R�!�4��0c�0�#�N[VDS�D0�;F!LwALO��CTO��kNN��M�OLR��END4�Lr+FVRC�ȺO�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�j�|������� ��������0B Tfx����� ��,>Pb t������� //(/:/L/^/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p����������ʿܿ� ���STD�LANG(�#�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9Kp]o��RBT'�OPTN�����
+DPN&�"/4/F/X/j/|/���/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/�? ?2?D?V?h?z?  ��?�?�?�?�?�?��=99E�$F�EAT_ADD �?	���/A~7@  	�8 @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n� �����������������""DDEMO �S/I   �8i_q��� ���
-7 d[m����� �/�/)/3/`/W/ i/�/�/�/�/�/�/? �/?%?/?\?S?e?�? �?�?�?�?�?�?�?O !O+OXOOOaO�O�O�O �O�O�O�O�O__'_ T_K_]_�_�_�_�_�_ �_�_�_�_o#oPoGo Yo�o}o�o�o�o�o�o �o�oLCU� y������� ��H�?�Q�~�u��� ����������� D�;�M�z�q������� ���ݟ�	��@�7� I�v�m��������� ٯ���<�3�E�r� i�{�������޿տ� ��8�/�A�n�e�w� �ϛϭ���������� 4�+�=�j�a�sߠߗ� �����������0�'� 9�f�]�o������ ��������,�#�5�b� Y�k������������� ����(1^Ug �������� $-ZQc�� ������ // )/V/M/_/�/�/�/�/ �/�/�/�/??%?R? I?[?�??�?�?�?�? �?�?OO!ONOEOWO �O{O�O�O�O�O�O�O ___J_A_S_�_w_ �_�_�_�_�_�_oo oFo=oOo|oso�o�o �o�o�o�oB 9Kxo���� �����>�5�G� t�k�}�������͏׏ ����:�1�C�p�g� y�������ɟӟ ��� 	�6�-�?�l�c�u��� ����ůϯ����2� )�;�h�_�q������� ��˿����.�%�7� d�[�mϚϑϣϽ��� ������*�!�3�`�W� iߖߍߟ߹������� ��&��/�\�S�e�� �����������"� �+�X�O�a������� ����������' TK]����� ���#PG Y�}����� �///L/C/U/�/ y/�/�/�/�/�/�/? 	??H???Q?~?u?�? �?�?�?�?�?OOO DO;OMOzOqO�O�O�O �O�O�O
___@_7_ I_v_m__�_�_�_�_ �_o�_o<o3oEoro io{o�o�o�o�o�o �o8/Anew �������� 4�+�=�j�a�s����� ď��͏����0�'� 9�f�]�o��������� ɟ�����,�#�5�b� Y�k���������ů� ���(��1�^�U�g� �������������� $��-�Z�Q�c�}χ� �ϫϽ������� �� )�V�M�_�y߃߰ߧ� ����������%�R� I�[�u������� ������!�N�E�W� q�{������������� JASmw ������ F=Ois�� ����///B/ 9/K/e/o/�/�/�/�/ �/�/?�/?>?5?G? a?k?�?�?�?�?�?�? O�?O:O1OCO]OgO �O�O�O�O�O�O _�O 	_6_-_?_Y_c_�_�_ �_�_�_�_�_�_o2o )o;oUo_o�o�o�o�o �o�o�o�o.%7 Q[���������*�!�M�  D�c�u����� ����Ϗ����)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9>K	  LQ gy������ �	-?Qcu �������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������������/APU Hk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S���$FEAT_D�EMOIN  VX�����X�k�_INDEXx�����k�ILECOM�P T��������f���S�ETUP2 U���Â�  �N �_AP2�BCK 1V��  �)T�"�1�%�U�X���C��� V����;�П_�ݟ� ��*���N�`��� ����I�ޯm����� 8�ǯ\��i���!��� E�ڿ�{�ϟ�4�F� տj����Ϡ�/���S� ��w���߭�B���f� x�ߜ�+�����a��� ���,��P���t�� ���9���]������ (���L�^������� ��G���k� ��6 ��Z��~��C ��y�2D� h����Q� u
//�@/�d/v/ /�/)/�/�/_/�/�/@?�/%?N?ȉ��P �� 2�*.V1RU?�?0*�?�?`
3�?�?�%�0PC�?|#O0FR6:O"ON�?sOKT���O �O8E�O�Lz�dO�O�&�*.F�?*_1	�:C_W\�O{_
[STM�_�_7B=@�_�]j_�_
[H�_2o�W� o�_�_�oZGIF �o�o�U�oaosoZJPG<�U(�o�o�JJS��0�Rs�j%
Ja�vaScript�CS�C��V0��� %Casc�ading St�yle Shee�tso�� 
ARGNAME.DT��
<�P\��p��q��󏟏�DISP	*��.ބ9���	��i�w�#�
TPEI?NS.XML��Ώ�:\��x�ځCus�tom Tool�bar��*�PAS�SWORDn��.FRS:\>���_��Password Config� �/ȯW�����4?"��� F�X��|������A� ֿe�������0Ͽ�T� �Mϊ�Ϯ�=����� s�ߗ�,�>���b��� ���'߼�K���o��� ��:���^�p��ߔ� #����Y���}���� ��H���l���e���1� ��U������� ��D V��z	�-?� c���.�R� v��;��q /�*/��`/��/ /}/�/I/�/m/?? �/8?�/\?n?�/�?!? �?E?W?�?{?O�?	O FO�?jO�?�O�O/O�O SO�O�O�O_�OB_�O �Ox__�_+_�_�_a_ �_�_o,o�_Po�_to �oo�o9o�o]ooo �o(�o!^�o� ��G�k ��� 6��Z�������� C����y����2�D� ӏh�������-�Q� �u������@�ϟ9� v����)���Я_��� ���*���N�ݯr�� ���7�̿[�ſϑ� &ϵ�J�\�뿀�Ϥ� ��E���i��ύϟ�4����$FILE_�DGBCK 1V���!���� < �)�
SUMMARY�.DG>���MD�:r߲���Di�ag Summa�ry����
CONSLOG�ߋߝ����6���Conso?le log7��	TPACCN,���%y����TP� Account�inX���FR6�:IPKDMP.'ZIP����
�;������Except�ion?����ME?MCHECK��������J�Memory Data����3l�)	F�TP)������L�mment T�BDG�L >I�)ETHERNET<�΁�����Etherne�t N�figur�a^���1DCSV�RF;!3L���% veri?fy allO��M.cDIF�FD*<���%=fdiff��|��CHG01����V/a�~/�- )2L/3/E/�/�{/�/"3�/�/�/^?� �/�?6V�TRNDIAG.�LS�?;?M?�?��ޢ1 Ope� L�og ��nost�ic��:�)�VDEV�2DAT��?�?�?�?bVi�sADeviceOKIMG�21�AO�SO�O�#~DIma�g�OKUP/@E�S.O�OFRS:�\._o]��Upd�ates Lis�to_���@FLEXEVEN��O�O��_a�Q UIF� Evb	@�_  �,�t)
PS�RBWLD.CM�o��ZR6oq_K�P�S_ROBOWE�Lh�:GIGE�	Oo�_�o��Gi�gEXo�N�A��)�aHADO�W�o�o�o|��S�hadow Ch�anges���a�<rRCMERARtYk ����p�CFG Erro�r�@tail� �MA����pSGLIB�����rI� St� A-�>�o�)r�ZD�op��o����ZD@�ad��3� <rNOTI��������Notific8�3�(f�AG��� �����;���_�� ����$���H�ݯ�~� ���7�I�دm�����  ���ǿV��z��!� ��E�Կi�{�
ϟ�.� ����d��ψ�߬�*� S���w�ߛ߭�<��� `�����+��O�a� �߅���8����n� ���'�9���]���� ��"���F�����|� ��5��Bk��� ��T�x� C�gy�,� P���/�?/Q/ �u//�/�/:/�/^/ �/?�/)?�/M?�/Z? �??�?6?�?�?l?O �?%O7O�?[O�?O�O  O�ODO�OhO�O_�O 3_�OW_i_�O�__�_ �_R_�_v_oo�_Ao �_eo�_ro�o*o�oNo �o�o�o�o=O�o s��8�\� ��'��K��o��� ���4�ɏۏj����� #�5�ďY��}���� ��B�ןf������1� ��U�g���������� P��t�	����?�ί c�򯇿��(���L���󿂿Ϧ�;�M��$�FILE_FRS�PRT  ���1�����\�MDONLY� 1Vp�(� �
 �)MD:�_VDAEXTP.ZZZN��������6%NO �Back fil�e ��(�S�6) ܿ7���[�$�hߑ�ֿ ��D�����z���3� E���i��ߍ��.��� R���v������A��� e�w����*�����`� ����+��O��s ��8�\� �'�K]�����`�VISBC�K��x���*.V�D�/pFR:�\�ION\DA�TA\��p�Vision VD�./<v/�/��/ ��/_/�/?�/*?�/ N?`?�/�??�?7?I? �?m?OO�?8O�?\O �?mO�O!O�OEO�O�O {O_�O4_�O�Oj_�O �_�_[_�_S_�_w_�_ o�_Bo�_foxoo�o�+o�oOoao�oV�LU�I_CONFIG7 Wp��{� $ �c��{ p�Xj|����y@p|x�o��� � 2�B��e�w������� D��������+� O�a�s�������@�͟ ߟ���'���K�]� o�������<�ɯۯ� ���#���G�Y�k�}� ����8�ſ׿���� ϶�C�U�g�yϋϝ� 4���������	ߠ�� ?�Q�c�u߇�߽߫� ��������)�;�M� _�q��������� �����%�7�I�[�m� �������������� ��!3EWi{ ������� /ASe�v�� ���z//+/=/ O/a/��/�/�/�/�/ �/v/??'?9?K?]? �/�?�?�?�?�?�?r? �?O#O5OGOYO�?}O �O�O�O�O�OnO�O_ _1_C_U_�Oy_�_�_ �_�_X_�_�_	oo-o ?o�_couo�o�o�o�o To�o�o);�o _q����P� ���%�7��[�m� �������L�ُ��� �!�3�ƏW�i�{���(����A�͐x��ʓ��$FLUI_D�ATA X�������D��RESULT� 2Y��#� ��T�/wi�zard/gui�ded/step�s/Expert ٟZ�l�~�������Ư�د������C�ontinue �with G7�ance�W�i�{��� ����ÿտ����ϋ ˒-̑��<�0 �M�<�����6\��.�psϧ� ����������%�7� I�[�m�,�M��ߦ߸� ������ ��$�6�H�Z�l�~�\�N�`�r�>��torch���� ��*�<�N�`�r��� ������y����� &8J\n��������������wproc��HZl ~������� /��2/D/V/h/z/�/ �/�/�/�/�/�/
?? ��7?{���@��TimeUS/DST&?�?�?�?�?�?�OO,O>OPObO%�EnablE��O�O �O�O�O�O__&_8_(J_\_n_˒8�F?0�_j?|?�624�?�_ o"o4oFoXojo|o�o �o�oqO�O�o�o 0BTfx��� �_�_�_�_w�-�?�?Region�R� d�v���������Џ����!�America<@�R�d�v� ��������П����!��qy��P��$��2Edi������� ʯܯ� ��$�6�H��Z�+ Touch Panel ��� (recommen��)h�����ѿ �����+�=�O�a� ��0�B���f�x��2acces/���� �/�A�S�e�w߉ߛ����,Conne�ct to Network����� �)�;�M�_�q���(���$���p�Ϛ����\!�ϐ0Int?roduct>�Q� c�u������������� �� /);M_q ������� 0?��0
��R #������� //(/:/L/^/�/ �/�/�/�/�/�/ ?? $?6?H?Z?�x3P:H�?l�?�?�? OO+O=OOOaOsO�O �O�Oh/�O�O�O__ '_9_K_]_o_�_�_�_ �_v?�?�?�_�?#o5o GoYoko}o�o�o�o�o �o�o�o�O1CU gy������ �	��_*��_N�ou� ��������Ϗ��� �)�;�M�_�p����� ����˟ݟ���%� 7�I�[��|�>���b� ǯٯ����!�3�E� W�i�{�������p�տ �����/�A�S�e� wωϛϭ�l��ϐ��� ����+�=�O�a�s߅� �ߩ߻��������¿ '�9�K�]�o���� ����������� ��� D�V��}��������� ������1CU �y������ �	-?Q�Z� 4�~�j����/ /)/;/M/_/q/�/�/ �/f�/�/�/??%? 7?I?[?m??�?�?b ���?�?�!O3OEO WOiO{O�O�O�O�O�O �O�O�/_/_A_S_e_ w_�_�_�_�_�_�_�_ �?�?�?�?LoOso�o �o�o�o�o�o�o '9K
_o��� ������#�5� G�Y�o*o<o��`oŏ ׏�����1�C�U� g�y�����\��ӟ� ��	��-�?�Q�c�u� ������j�|���𯲏 �)�;�M�_�q����� ����˿ݿ￮� �%� 7�I�[�m�ϑϣϵ� �������ϼ���B� �i�{ߍߟ߱����� ������/�A�S�d� w����������� ��+�=�O��p�2� ��V߻������� '9K]o��� d�����#5 GYk}��`�� ������/1/C/U/ g/y/�/�/�/�/�/�/ �/�?-???Q?c?u? �?�?�?�?�?�?�?� O�8OJO?qO�O�O �O�O�O�O�O__%_ 7_I_?m__�_�_�_ �_�_�_�_o!o3oEo ONO(Oro�o^O�o�o �o�o/ASe w��Z_���� ��+�=�O�a�s��� ��Vo�ozoďo� '�9�K�]�o������� ��ɟ۟ퟬ�#�5� G�Y�k�}�������ů ׯ鯨���̏ޏ@�� g�y���������ӿ� ��	��-�?���c�u� �ϙϫϽ�������� �)�;�M���0��� T�����������%� 7�I�[�m���Pϵ� ���������!�3�E� W�i�{�����^�p߂� ����/ASe w�������� �+=Oas� ��������/ ��6/��]/o/�/�/�/ �/�/�/�/�/?#?5? G?X/k?}?�?�?�?�? �?�?�?OO1OCO/ dO&/�OJ/�O�O�O�O �O	__-_?_Q_c_u_ �_�_X?�_�_�_�_o o)o;oMo_oqo�o�o TO�oxO�o�O�o% 7I[m��� ����_�!�3�E� W�i�{�������ÏՏ 珦o��o,�>��e� w���������џ��� ��+�=��a�s��� ������ͯ߯��� '�9���B��f���R� ��ɿۿ����#�5� G�Y�k�}Ϗ�N����� ��������1�C�U� g�yߋ�J���n����� ��	��-�?�Q�c�u� ����������� �)�;�M�_�q����� ���������߮����� 4��[m��� ����!3�� Wi{����� ��////A/  $�/H�/�/�/�/�/ ??+?=?O?a?s?�? D�?�?�?�?�?OO 'O9OKO]OoO�O�OR/ d/v/�O�/�O_#_5_ G_Y_k_}_�_�_�_�_ �_�?�_oo1oCoUo goyo�o�o�o�o�o�o �O�O*�OQcu �������� �)�;�L_�q����� ����ˏݏ���%� 7��oX�|�>���� ǟٟ����!�3�E� W�i�{���L���ïկ �����/�A�S�e� w���H���l�ο���� ��+�=�O�a�sυ� �ϩϻ����Ϟ��� '�9�K�]�o߁ߓߥ� �����ߚ��߾� �2� ��Y�k�}������ ��������1���U� g�y������������� ��	-��6��Z �F����� );M_q�B� �����//%/ 7/I/[/m//>�b �/�/��/?!?3?E? W?i?{?�?�?�?�?�? ��?OO/OAOSOeO wO�O�O�O�O�O�/�/ �/�/(_�/O_a_s_�_ �_�_�_�_�_�_oo 'o�?Ko]ooo�o�o�o �o�o�o�o�o#5 �O__z<_��� �����1�C�U� g�y�8o������ӏ� ��	��-�?�Q�c�u� ��FXj̟��� �)�;�M�_�q����� ����˯��ܯ��%� 7�I�[�m�������� ǿٿ���������E� W�i�{ύϟϱ����� ������/�@�S�e� w߉ߛ߭߿������� ��+��L��p�2� ������������ '�9�K�]�o���@ߥ� ����������#5 GYk}<�`�� ���1CU gy������� �	//-/?/Q/c/u/ �/�/�/�/�/��/� ?&?�M?_?q?�?�? �?�?�?�?�?OO%O �IO[OmOO�O�O�O �O�O�O�O_!_�/*? ?N_x_:?�_�_�_�_ �_�_oo/oAoSoeo wo6O�o�o�o�o�o�o +=Oas2_ |_V_���_��� '�9�K�]�o������� ��ɏ�o����#�5� G�Y�k�}�������ş ������C�U� g�y���������ӯ� ��	��ڏ?�Q�c�u� ��������Ͽ��� �)�����n�0��� �Ϲ���������%� 7�I�[�m�,��ߣߵ� ���������!�3�E� W�i�{�:�L�^���� ������/�A�S�e� w���������~����� +=Oas� ��������� ��9K]o��� �����/#/4 G/Y/k/}/�/�/�/�/ �/�/�/??�@? d?&�?�?�?�?�?�? �?	OO-O?OQOcOuO 4/�O�O�O�O�O�O_ _)_;_M___q_0?�_ T?�_x?z_�_oo%o 7oIo[omoo�o�o�o �o�O�o�o!3E Wi{�����_ ��_���oA�S�e� w���������я��� ���o=�O�a�s��� ������͟ߟ��� ���B�l�.����� ��ɯۯ����#�5� G�Y�k�*�������ſ ׿�����1�C�U� g�&�p�J��Ͼπ��� ��	��-�?�Q�c�u� �ߙ߽߫�|������ �)�;�M�_�q��� ���xϊϜϮ���� 7�I�[�m�������� ����������3E Wi{����� ������ �b $�������� //+/=/O/a/ �/ �/�/�/�/�/�/?? '?9?K?]?o?.@R �?v�?�?�?O#O5O GOYOkO}O�O�O�Or/ �O�O�O__1_C_U_ g_y_�_�_�_�_�?�_ �?o�?-o?oQocouo �o�o�o�o�o�o�o (o;M_q�� ��������_ 4��_X�o������� Ǐُ����!�3�E� W�i�(������ß՟ �����/�A�S�e� $���H���l�n���� ��+�=�O�a�s��� ������z�߿��� '�9�K�]�oρϓϥ� ��v��Ϛ����ҿ5� G�Y�k�}ߏߡ߳��� �������̿1�C�U� g�y���������� ��	������6�`�"� �������������� );M_�� �����% 7I[�d�>��� t����/!/3/E/ W/i/{/�/�/�/p�/ �/�/??/?A?S?e? w?�?�?�?l~�� O�+O=OOOaOsO�O �O�O�O�O�O�O_�/ '_9_K_]_o_�_�_�_ �_�_�_�_�_o�?�? �?VoO}o�o�o�o�o �o�o�o1CU _y������ �	��-�?�Q�c�"o 4oFo��joϏ��� �)�;�M�_�q����� ��f��ݟ���%� 7�I�[�m�������� t�֯������!�3�E� W�i�{�������ÿտ �����/�A�S�e� wωϛϭϿ������� �Ư(��L��s߅� �ߩ߻��������� '�9�K�]�ρ��� �����������#�5� G�Y��z�<ߞ�`�b� ������1CU gy���n��� �	-?Qcu ���j�����/ �)/;/M/_/q/�/�/ �/�/�/�/�/?�%? 7?I?[?m??�?�?�? �?�?�?�?�/�*O TO/{O�O�O�O�O�O �O�O__/_A_S_? w_�_�_�_�_�_�_�_ oo+o=oOoOXO2O |o�ohO�o�o�o '9K]o��� d_�����#�5� G�Y�k�}�����`oro �o�o���o�1�C�U� g�y���������ӟ� ����-�?�Q�c�u� ��������ϯ��� ď֏�J��q����� ����˿ݿ���%� 7�I��m�ϑϣϵ� ���������!�3�E� W��(�:���^����� ������/�A�S�e� w���ZϬ������� ��+�=�O�a�s��� ����h��������� '9K]o��� �����#5 GYk}���� �����/��@/ g/y/�/�/�/�/�/�/ �/	??-???Q?u? �?�?�?�?�?�?�?O O)O;OMO/nO0/�O T/VO�O�O�O__%_ 7_I_[_m__�_�_b? �_�_�_�_o!o3oEo Woio{o�o�o^O�o�O �o�o�_/ASe w������� �_�+�=�O�a�s��� ������͏ߏ�o�o �o�H�
o������� ��ɟ۟����#�5� G��k�}�������ů ׯ�����1�C�� L�&�p���\���ӿ� ��	��-�?�Q�c�u� �ϙ�X���������� �)�;�M�_�q߃ߕ� T�f�x����߮��%� 7�I�[�m����� ��������!�3�E� W�i�{����������� ����������> �e w������� +=��as� ������// '/9/K/
.�/R �/�/�/�/�/?#?5? G?Y?k?}?�?N�?�? �?�?�?OO1OCOUO gOyO�O�O\/�O�/�O �/	__-_?_Q_c_u_ �_�_�_�_�_�_�__ o)o;oMo_oqo�o�o �o�o�o�o�o�O�O 4�O[m��� �����!�3�E� oi�{�������ÏՏ �����/�A� b� $��HJ���џ��� ��+�=�O�a�s��� ��V���ͯ߯��� '�9�K�]�o�����R� ��v�ؿ꿮��#�5� G�Y�k�}Ϗϡϳ��� ���Ϩ���1�C�U� g�yߋߝ߯������� ���ȿ�<���c�u� ������������ �)�;���_�q����� ����������% 7��@��d�P� ����!3E Wi{�L���� ��////A/S/e/ w/�/HZl~�/� ??+?=?O?a?s?�? �?�?�?�?�?�OO 'O9OKO]OoO�O�O�O �O�O�O�O�/�/�/2_ �/Y_k_}_�_�_�_�_ �_�_�_oo1o�?Uo goyo�o�o�o�o�o�o �o	-?�O_"_ �F_������ �)�;�M�_�q���Bo ����ˏݏ���%� 7�I�[�m����P�� t֟����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ㿢� �Ɵ(��O�a�sυ� �ϩϻ��������� '�9���]�o߁ߓߥ� �����������#�5� ��V��z�<�>���� ��������1�C�U� g�y���J߯������� ��	-?Qcu �F�j����� );M_q�� ������//%/ 7/I/[/m//�/�/�/ �/�/���?0?� W?i?{?�?�?�?�?�? �?�?OO/O�SOeO wO�O�O�O�O�O�O�O __+_�/4??X_�_ D?�_�_�_�_�_oo 'o9oKo]ooo�o@O�o �o�o�o�o�o#5 GYk}<_N_`_r_ ��_���1�C�U� g�y���������ӏ�o ��	��-�?�Q�c�u� ��������ϟ០� �&��M�_�q����� ����˯ݯ���%� �I�[�m�������� ǿٿ����!�3�� ��x�:��ϱ����� ������/�A�S�e� w�6��߭߿������� ��+�=�O�a�s�� DϦ�h�������� '�9�K�]�o������� ����������#5 GYk}���� ��������CU gy������ �	//-/��Q/c/u/ �/�/�/�/�/�/�/? ?)?�J?n?02? �?�?�?�?�?OO%O 7OIO[OmOO>/�O�O �O�O�O�O_!_3_E_ W_i_{_:?�_^?�_�_ �O�_oo/oAoSoeo wo�o�o�o�o�o�O�o +=Oas� �����_�_�_� $��_K�]�o������� ��ɏۏ����#��o G�Y�k�}�������ş ן������(�� L�v�8�������ӯ� ��	��-�?�Q�c�u� 4�������Ͽ��� �)�;�M�_�q�0�B� T�f��ϊ�����%� 7�I�[�m�ߑߣߵ� �߆������!�3�E� W�i�{�������� �Ϧϸ����A�S�e� w��������������� ��=Oas� ������ '����
�l.��� �����/#/5/ G/Y/k/*|/�/�/�/ �/�/�/??1?C?U? g?y?8�?\�?��? �?	OO-O?OQOcOuO �O�O�O�O�O�?�O_ _)_;_M___q_�_�_ �_�_�_�?�_�?o�? 7oIo[omoo�o�o�o �o�o�o�o!�OE Wi{����� �����_>� ob� $o&�������я��� ��+�=�O�a�s�2 ������͟ߟ��� '�9�K�]�o�.���R� ��Ư������#�5� G�Y�k�}�������ſ �������1�C�U� g�yϋϝϯ��π�ʯ �����گ?�Q�c�u� �ߙ߽߫�������� �ֿ;�M�_�q��� ������������� ���@�j�,ߑ����� ��������!3E Wi(����� ��/ASe $�6�H�Z��~��� //+/=/O/a/s/�/ �/�/�/z�/�/?? '?9?K?]?o?�?�?�?��?�?���OE��$FMR2_GR�P 1ZE�� �C4�  B�� 	 �� VOhLS@F@ ~EE���B~A�:�{A�L�FZ!�D�`�D�� �BT��@����M?�  �O�<S@�6����B���5�Zf5�ES<Q�MA�  _0[�BHT�@JQ@�3�3@�TPXS�<RDx_�]S@@OQ�_�N��_�_RA<�z�<��ڔ=7�<��
;;�*�<����M8ۧ��9k'V8���8���7ג	8(���_?o�_<o�uo`o�o�o�o�',B_�CFG [9KT�hB�o/�iNO� 9J
F0�cq hp�lRM_C�HKTYP  �)A� A@C@�0+ARO=M~p_MIN�p�#W���p�oPX,@�SSB�c\E TF��%��s���eTP_D�EF_OW  ��$AC$�IRCO�M�p5��$GENOVRD_DO�v��!b�THR�v �d�dh�_ENB�T� h�RAVC�2C]�w�p �@vE� ��o$��L2��C�fZ �ȁOU*5@c9LkqfH9�fE<�p�O��d��ԟ��#C�  AD+�1���L�\�@OAC�B�gAI�iI���.ɀSMT2Cd։E@��p'��$HOST�C�b1e9I�pй�/R@ MC�$�?����&  �27.0M�16�  e-�z������� ��h�����:�ѿ�˳	anonymous>�l�~ϐϢ� ���"��Q@����+� -��a�B�T�f�xߊ� Ϳ��������ߡ�K� ,�>�P�b�t������ �������5��(�:� L��	����������� ��� $6H�� ����������� � c�DVhz ���������
/ /_q���m/� �/�/�/�/�/7?*? <?N?`?�/���?�? �?�?�?3/E/W/i/k? \O�/�O�O�O�O�O? �O�O_"_4_WO�?N_ |_�_�_�_�_OO+O �_?_0osOTofoxo�o �o�O�o�o�o�oo ]_>Pbt���_ �_�_��Go(�:� L�^��o��������ʏ �o�1�$�6�H�Z����ߡENT 1f~��  P!�.��  ����֟ ş������B��N� )�w���_�����䯧� �˯,���b�%��� I���m�ο�����ǿ (��L��p�3�iϦ� ���ύ��ϱ����� ��G�l�/ߐ�Sߴ�w� �ߛ��߿���2���V���z�=�QUIC�C0��c�u����1 �����&���2'����v�!ROUT�ERw�S�e���!�PCJOG�����!192.16?8.0.10���?CAMPRT���!1 >%R�T��BT� !�Software� Operator Panel��{�NAME �!��!ROB�O0S_CFG� 1e�� ��Auto-started�t/FTP��� ޏ����/#/5/ ~�Y/k/}/�/��/F/ �/�/�/??1?�pw ��|?�/��?�?�? �?�?�/O0OBOTOfO �?O�O�O�O�O�O�O ����qOG_�?�_ �_�_�_�_�O�_oo (o:o]_�_po�o�o�o �o�o__1_C_Eo6 y_Zl~��eo� ����1�D�V� h�z������o�o�� �
�M.�@�R�d�v� 9�������П����� �*�<�N�`�r���Ǐ ُ���ޯ!���&� 8���\�n�������ǯ I�ÿ����"�4�w� ��������������� �����Ͽ0�B�T�f� xߛ�߮��������� �K�]�oρσ�t�� ����������� (�:�L�o��������������_ERR� g&����PDUSIZ  q�^���>$W�RD ?eR���  guestq�dv�����SCD_GROUP 3he� i{�IFT�$PAOMP� _SHvEDS $C�COM��TTP_AUTH 1i� <!iPendan���q��n1!KARE�L:*���K�C//'/�VI�SION SET� �/\/m6!�/�/�/ ��/�/�/�/7?? ?�m?D?V>�CTRL� j�8q�
�q�FFF9E�3y?P�FRS:DEFAULT�<�FANUC �Web Server�:�2R�L^ �<YOkO}O�O�O�O���WR_CONFI�G k��?�?��IDL_�CPU_PC@�q�B�S�%P BH�UMIN\�)UGNR_IO��2q��	PNPT_SI�M_DO[Ve[S�TAL_SCRN�[V ��6oQTPM?ODNTOL�We[>ARTY|X%QjVy .�ENB�W�
SOLNK 1l -o?oQocouo�o|�obMASTEZP�ijUOSLAV�E m�eRA?MCACHE�o�R}O�O_CFG�o�csUO� rCMT_OP@]R
�OsYCL�o+u�0_?ASG 1n�G>
 �o���� ��*�<�N�`�r���p�����k�rNUM15	
rIP�owRTRY_CNZ<+u�Q_UPD1,a�� r8pro��n� g�� PRCA_ACC 2p��  Wk) �(C�  �� 5
� 6�q��,�Rᛖ3� G)������ ˝�}�BUF001 �2q�= h/�u0  u0h@��O�`�o�������������������iU~�~�!~�1~�UB~�Q~�b~�r~�U�~��~��~��~�U�~��~��~����j����,u0�(sjS��u�u0/�Exj�������������ƪ����������k�f�)u0K�)�@k8n�@l��f��f͆��j��톴��g��U��.��=��N���]��n��}� ]8S�8h� ���2���$�)�-� )�5�)�=�)�E�)�M� )�U�)�]�)�e�)�m� )�u�)�}������ �����¥��­� �µ��½���Š��͠���ՠ��ݠR�"��!�SX졉��� ������	��	���N0' �s�h,�	�5�	�=�	�E� 	�M�	�U�	�]�	�e��tp �l��t�t�� �|�n�   ������ҕ��ҝ��� ������ҵ��ҽ��� Ű��Ͱ��հ��ݰ�� �)�����)������3��+�2�-�;� 2�=�K�2�M�[�2�]� k�2�m�{�2�}��Ò� ���Ò❢�Ò⭢�� �⽢�Ò�͢�Ò�ݢ ��墋���Ò���� ������%�� -�;��=�K��M�[� �]�k�\l�{�z�}� \���Ӓ򕲣Ӓ� �Ӻ��Ӻ�Ų�Ӻ� ղ�Ӻ����2�����	T��q2r� Q4�<�5\\<\�PS]R}�HIS��t� ܛ�� 2023-08�-16\+g7�\;�����Zh2\:{��0: b�*<N�W�� ��7���������R	AS �	A� ��P/#/|=3,k�} j/|/�/�/�/�/�/�/ �/?C/U/B?T?f?x? �?�?�?�?�?�??-? O,O>OPObOtO�O�O �O�O�?O�O__(_ :_L_^_p_�_�_�O�O �O�_�_ oo$o6oHo Zolo��k�w�w� �d{o�o�o�U9: c��9` K]o]ox�� ����Sd �b 	 !��G��_�_��� ����ŏ׏����� 1�h�z�g�y������� ��ӟ���	�@�R�?� Q�c�u���������ϯ ��*��)�;�M�_� q������������ ��%�7�I�[�m�� ��o�e��o�o��  C	��)�;�C=�l�~ߐ�~�� ������� ����" ��	 ��g�y�׿鿯� ��������	��-�?� Q������������� ����)`�r�_ q������� 8J\I[m ������"4 !/3/E/W/i/{/�/�/��/�/�eI_CFG� 2u�� H�
Cycle T�ime�Bus=y�Idl2��min�+R��Up�&�Re�ad7Dow�+8'?6p<1�#Co�unt�	Num� �"����<���1�aPROG�"-v������?�?�O!O3OEOWO29�eS�DT_ISOLC�  ���Y�Z���$J23_DSP_ENB  �K�PЫ@INC w��M�Ә@A   ?��=���<#��
�A�I:�o  �A_(_��_P_�G�0�GROUP 1xv�K!�< P�C��_X_?��?�_��Q�_o!o3o�_ Woio{o�o�@_b[�IN_AUTO � ���J�@POS�REC�C�b71�hK�ANJI_MAS�K�f�jKAREL?MON y�˰?��yRok}���(�.)r�3z�7�C����u�ouCL_L��`NUM�@
��@K�EYLOGGIN�G�`����Q�E�0L�ANGUAGE ���q���DEFAULT l���LG�!{�:�72��x�@� � 8P�H  �V��'0���Л��ycOU�;��
�(UT1:\�� ��.�@�W��d�v����������(�Z���LN_DISP |�O48�_|�_!�OCTOL`����Dz�0�A�Av�GBOOK }���dޔR��ᑮ�X ٌү�����,�<�0��P�N�*�	��ۉ��QmK��aO�A��_B�UFF 2~�K ���235ݿ�� R���17�'�T�K�]� �ρϓ��Ϸ������� ���#�P�G�Y߆��C~��DCS ��9 �B�AK�����%�� ���$��IO 2���� !Z�Q�]�m������� �������!�5�E�W� i�}����������������8�ER_ITM�Nd�ofx�� �����, >Pbt����8�p�;SEV�`�M]7TYP�NU�6/H/Z/��aRST�(���SCRN_F�L 2�F��0� ���/�/�/??(?:?Fk/TP>��O%"M=NGNAM�Dǥq�n��UPS)�GI� �	��E�1_LO�ADPROG �%g:%	T_AR�CWELDG?�MAXUALRM%�,�a���E
B�1'_PR�4�` ��L�@C,����hO����%��ODoPP 2�.�� �ؖ	%/�O �O�O�O_-__Q_<_ u_X_j_�_�_�_�_�_ o�_)ooMo0oBo�o no�o�o�o�o�o�o %[Fj� �������3� �W�B�{���p����� Տ��ʏ���/��S� e�H���t�������� Ο��+�=� �a�L� ��h�z�����߯ʯ�����9�$�]�HDBGDEF �YE���eOu�_LDXD�ISA�0f;6�ME�MO_AP�0E {?g;
 �� F������/�A�S��e�@FRQ_CF�G �YG��AM F�@���H�<�ԃd%h���yϋ��B��YKL��*�/� **: (�H��-���H�S�e� �߉ߛ��߿�����J� YE'� �N�<�R�`�,(�ߥ������ �����*��N�5�r� ��k�����������~JISC 1�g9� �P�JL���`�K���� _M?STR ����SCD 1�ֽ� �/�S>wb� ������// =/(/M/s/^/�/�/�/ �/�/�/?�/ ?9?$? ]?H?�?l?�?�?�?�? �?�?�?#OOGO2OkO VOhO�O�O�O�O�O�O _�O_C_._g_R_�_ v_�_�_�_�_�_	o�_ -ooQo<ouo`o�o�o �o�o�o�o�o;��MJPT��1���i�{�w^sMI�R 1����p ��L���.s< ��?O��.q?y3�\�N��  ����P���.���©� &��5C��o.q���~ �+yH��@�b���v� ��Ə珺����ҏ D�b�4�^���b����� П��؟�+y����L� ^�����g�q���ͯ k�ů�����K�-� ~�����5�W�ɿ���� ׿ϯ��G�-�?�a� c�q�����g�yϛ�� ����U�;�]ߋ�q� ���ߣϵ���߽� ?���3�=��a��� ����������J�\� �����e�w����i� ��������I+�| ��3U����� �E+=_��o^pKdq�j{ � �\rLTARkM_��ju�p��xtop/$^pME�TPU  .r��]qNDSP?_ADCOL3%��>.CMNTT/ �G%FNp t/E'FS�TLI�/�'MST ���/xs� ?|
4G%POSCF�'=.PRPMs/9[STR 1�j}4�q<#�
�16q�5�? �7�?�?�?�?�?�?�? .OO"OdOFOXO�O|O��O�O�O�O_�AG!S�ING_CHK � �/$MODAQ��jy��@U�DEV 	jz	�MC:t\HSI�ZE3 ��@UTA�SK %jz%$�12345678�9 �_�U>WTRI�fp�j{ lju% �8oh+oloOm�t�S�YP�Q{uVT?SE�M_INF 1���XQ`)AT&FV0E0uo��m)�aE0V1�&A3&B1&D�2&S0&C1S�0=�m)ATZ�o@'tHDl�a`o�#xA������ �oC��o ,��P������� �֏?�Q�8�u�(�:� ��^�p��������)� `�M�����>����� ˯ݯ�����Ɵ؟� [���������h�ٿ �������3����i� �.�@�����v���� ���пA���e�L߉� ��NϿ�rτϖϨ�� ��=�O��s�&ߗ�R��������m_NIT�OR� G ?�[ �  	EXESC1�"3�2:�3:�E4:�5:�`<�7:�8:�9:�5�ҟ� 9��E��Q��]�� i��u������T���2��2��2��U2��2��2��2��U2��223���3��3E�@QR_G�RP_SV 1���k (�A?�=��!4 �{ ����Q_D��^�IO/N_DBJP�N]�!_  �@�cX�? /� ��O��@�cX��N ]��]GOQ�hT-ud1�U����a�PL_NAME �!e��!�Default �Personal�ity (fro�m FD)�R�R2� 1�L?�XL�x�hP d�"J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�?�?�?�?aS2F/�?O O%O7OIO[OmOO�OaR<�?�O�O�O�O_ _'_9_K_]_o_�_�%�F�O�^
�_�_�P�_oo/oAoSo eowo�o�o�o�o�o�o �o�_�_Oas �������� �'�9�K�]�,>�� ����ɏۏ����#� 5�G�Y�k�}�������� H�6 H?�b H\��� �  �����d ܓĐ�#��E�S�Ő ���=����������� ��ٯϯ�� ��5�W�� z������	`ï��Ͽ|ῠ�:�oA!"���%�7� A'�  Lɨ�'tw�.�������e~� �G��hȟ���ϰ���@�����
�C��R�� 1��u��?@ � ���~�� @D�  ��?��Ӂ�?�����A��6Ez  x�ј��;�	l���	 �@�� 0�vw�� ���� � � ���� J��K ���J˷�J� ��J�4�JR��<(�7'��d�� @��S�@�;fA�6A��A1UA��X@��O��=�N��f������T;�f��X����E��*  ���  �5��>������ҘM�� �?���#�������6�w�(�� �>�=���P�H�Y�u�u�(y��u��Ï�5߫�N�	'� � ���I� �  ��Y�L�:�È~��È=���~Q��� <���� � ?� �e���?����I�p�~ėe��z��@!�p@�a�@��@��@��C��C�� �� ��B��Cz��d�@�7������3���� K�L�����I�@�m�D�՚��������(
%Y:�a�  =�x?��ffd�K/]/� !���/�+R�8Y �/�*>��=��I� ���&��6)�����Ԟ_>���A!E�<�2�!<"7�<�L��<`N<D��<��,-�j?y/�����"I��?fff?m?&��0q�@T싹1?��`?Uȩ?X��1W	�1�� ����?��O�7��|/ QO<OuO`O�O�O�O�O��O�O�O_W�5F � _S__w_�?�_I�j_�_fXHmN H�[�YG� F���_oo
oCo.o goRo�ovo�o�o�o�o �et}�o`��_T�_ {�o����t?� ��/��S�>�w�b�AU��Uɲ�Cq� ֏m���������XD�/�W	ç��®�V��BH� �� T���� ������@I��Y�@n�@���@: @l��?٧]��� ��%�n��߱���?=�=D��������@�oA��&{C/� @�U���+J8���
H��>���=3H��_�E� F�6�G���E�A5F�ĮE��m�����fG���E��+E���EX����>\��G�ZE�M��F�lD�
 �п���
���.��R� =�v�a�������п�� ��߿��<�'�L�r� ]ϖρϺϥ������ ����8�#�\�G߀�k� �ߏߴ���������"� �F�1�j�U�g��� �����������B� -�f�Q���u������� ������,P; t_������ �:%7p+�=(-�4�t-1����]3�ϩx����4 �{�<����0+#����jb/+/1E�䴛|�0G+E)��/s/�/�/�/�,.uPe2P�.q(?{@4?^?I?�?m9F ��?��?�?�?�?�?�?��$ OOLO7OpO[O�O;? �O�O�O�Le�O�O�1__A_g_U_1) m__�_�_�_�_�_j�  2 H�6f��H�@",c\���1B������Bȓ���A��@��so��w��o �o�o�o�o1v#o5o�,>P`|��J�T�����Aotc��
 `�� ����&�8�J�\��n�������#�rr����H-��$M�R_CABLE �2��( TV`2T0aa@3 a?w��ab��{��?`B?`C �3!OM��`B���nr���+�r3 E�V�3&���J`�N`By�S`�O
�v7���E!��Ņt E��A%W�i�Z`��J`CW`9-���7�򏒞OF��$0�����*!��:�B:�C�/�7u 7�����RouD�\,������Z� +u�M�_�į��ͯ�� ���ݯ�T�O�%�q�@I�[����ɿ7� �!���(�:�1(�iϸ{ύ�1(*��*�* ݃OM �����HN�'��l%% 2345?678901���Ł ����3 :�ba�3 3!
כ��not sent� ��?�W�%�TESTFECS7ALG>�eg0*ba�d�ԈqF�F�F�0�0k~h������1(9UD1:\�maintena�nces.xml��_�  �z��DEFAULT��l݂GRP 2���  p�tg3%�  �%1st� mechani�cal chec�k�3!�������U� �j7�I��[�m��3"��controller���������T(���0!3E��M��m3""8�3 ���U�������P
C��3�W����������C���ge��. battery�G/�U	tI/[/m//�/���Supply? greasQ�/����#<��!�/�U8/??1?C?U?z���cabl�/�/�?,(
�/�?�?�? OO�����?�?��?�O�O�O�O�O%@A$�O_Ը׿4_ �O Y_k_}_�_�_�O�__ &_8_�_o1oCoUogo �_�o�_�_�_�o�o�o 	jo�oQ�o@�o �����0�� f;��_�q������� �ˏ�,��P�%�7� I�[�m��������ǟ �����!�3���W� ������ܟ��ïկ� ��H��l�~�S���w� ����������2�D� �h�=�O�a�sυ�Կ ����
������'� 9�Kߚ�o߾����Ϸ� ��������N߶�5�� $��}������� ����J��n�C�U�g� y�����������4� 	-?Q��u�� �������� f;��q��� ���,/Pb7/ �[/m//�/�/��/ /(/�/L/!?3?E?W? i?�/�?�/�/ ?�?�? �?OO/O~?SO�?�? �?�O�O�O�O�O2O�O _hO_�Oa_s_�_�_ �_�O�_�_._oR_'o 9oKo]ooo�_�o�_�_ �oo�o�o#5�l�b	 TCp�� �o������!� 3�E�W�i�{������� ÏՏ�����/�A� S�e�w���������џ������+�=� � ��a?�  @�a �x�������fd�ɯۯ�h*�** �a�f�� ?�A�S�e�'������������o�c$�¿ �"�4���X�j�|�ƿ ؿ�P�������D�� 0�B�Tߞϰ�ߜ߮� ��
ߔ�����d�v� ��&�t���Z�������*�<�j�$MR�_HIST 2���e;�� 
 \��b$ 2345678901K�S��
�J�9�o����s� ���o(����^ p�9K����  �$6�Z~ �G�k���/ �2/D/�h//�/�/�U/�/ �SKCFM�AP  �eU>���z z ��/�%ONREL  z$;��!� �"EXCFENB%7q
�#�%>1FNCE?�74JOGOVLI�M%7d;�0�"KE�Y%7�5�5_P�AN$8�2�2�"RU�N�<�;SFSP�DTYPe805�#S�IGN%?74T1M�OT�?41�"_C�E_GRP 1��e�#C�[p���O z#|O�O&D�O�O�O_ _�O>_�ON_t_+_�_ O_�_�_�_�_o�_(o �_Lo^oEo�o9o�o�o �o�o�o�o�o6�k��!QZ_EDIT�"D�'CTCOM_�CFG 1��-�H5��� 
vq_/ARC_B2%Ep9�T_MN_MOD�E"F�P9UAP�_CPL�T4NO�CHECK ?^�+ �/ S� e�w���������я� ����+�=�O�a�;�NO_WAIT_�L!GkwV@NT~qѩ�+�ez#��_E�RR`A2��)�!� ��
��.���1S�e�Ԏ��pOᓫ�| �(C�+qC�B�F���=�B[~�W<=/�!}Zx)<�0�� ?�k�Яk�0���ڒPARAM⒬�+�O�,S�>�8�!p��� = ���� ������ۿ�ɿ��#��5��Y�k�G�=����ϯ�B���BODR�DSP�s$FP8OF�FSET_CAR8ap$�	�DIS��wS_A�pARK"G�lyOPEN_FI�LE5�$A�qlv�pO�PTION_IO��?�1��M_PRGw %�*%$*��l��i�WOU��fGP���	�z$��G   2P�#���#�	 �x(#��z#����RG_DS�BL  3��!�̚����RIENTkTO$0z!C�0��!A ��UT_S/IM_D���"P����V��LCT ����hr�q�z%d��_PEX �8�+��RAT � dP5|+��UP ���|��������z T��z z 2�1֡��$�2_C�L�XL�x��%���+= Oas����� ��'9K]o�z'2��� ��
//./@/R/ã �|/�/�/�/�/�/�/��/??0?B?�il&@k/|>��|?�?ϒP�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �?�?_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo�O�OTofoxo�o �o�o�o�o�o�o�,>Pb��Co=�!���}!�����~ ����}�}��W�B�{�.�$�p������� ��ҏ؏���n���<�K�I�p�	`��~���<����:�o�����ҟ���o�A� � �i�'��.��Z��a��e?b[ ������� e���q��������˯��������Os�1�� �� � ���l�@ ��]��G� @D� M Z�?�`�F�?���b���D�  Ez�|�Y5�  ;�	�lr�	 ��@� c0g�h��� �V��� � � ��в��H0#H���G�9G��ģG�	{Gkf���S��,̖��C��\�%�D�	� D@ D�	������  ?�5��>t�[��ù�b�tφ� B���Bp{�=!����O�^���8��� а������f��6���:�(:��:��]�T����p��	'� �� ��I� ��  ���=���Ͳ���^���� <��� �� � ��*�^��u�^��5���N��\�&���ht�?���C��C�����B[���J���i0�Z��@������������������
�@��2�v���_�\�G� ��k����������������:!���x?�ff%�"��C [�Wi��8��<�
>���n� ��IкX��������<��$�>���
��<2�!<"7��<L��<`N�<D��<��,0�/>`����
�?fff?2�?y&l��@T�~�?�`?Uȩ?Xǎ�9��g s���b��`��P�� A//:/%/^/I/�/ m/�/�/�/�/�/�/? �/6?���/?�?+8HmN H[���G� F���? �?�?�?O�?,OOPO ;OtO_OqO�O�E9��M �O%�S?_w?@_�Od_ v_�_�_9�_�_[_�_ �_oo<o'o���fb�wkC6o�o2o�o�m?���o�o	,�o��çs��sm��H����Z�d��`�a�q@I����@n�@���@: @l���?٧]j ���%�n��߱���=��=D�ɺ�p���@�oA�&�{C/� @��U� �+J8���
H��>���=3H��_�
� F�6�G���E�A5F�ĮE��2��D���fG���E��+E���EX�Z�D�>\��G�ZE�M��F�lD�
 [���iϏ���ޏ� �;�&�_�J�\����� ����ݟȟ���7� "�[�F��j�����ǯ ��į���!��E�0� i�T�y�����ÿ��� ҿ���/��,�e�P� ��tϭϘ��ϼ���� ��+��O�:�s�^ߗ� �ߔ��߸������ � 9�$�I�o�Z��~�� ������������5��r=(�q4�9�����j�"�3�ϩxZ�l��q4 �{��<���q�0+#����Φ�jb����1E�䴛|[
	�J8n\���EP*P��A�O�@�@�#G2 �M�T�x����r$ ��/�5/ /Y/  �O�/z/�/�,e�/�/��/�/?,??�A) 2?D?z?h?�?�?�?�:�  2 H�6f�vH��3\��v1Boacao`B�XpWpA�p@so8OJO\OnO�O�O�M�CP/�O�OP�O__%\�vN$%�p�p�A4T�3�u
 %__�_�_ �_�_�_�_�_o!o3o`EoWoio�z7R�����H-��$PA�RAM_MENU� ?
��  M�NUTOOLNU�M[1�w�`F��`�`�iAWE�PCR�`.$INCH_RATE�`�SHELL_C�FG.$JOB_�BASp W�VWPR.$CENTER_RIr��`$tAZIMUT�H OPTB�a�$tELEVATI_ON TC�a$t�DWqTYPE �SNqARCLI�NK_AT(pST�ATUS�c�y__�VALUq�`L�EP�a.$WP_ �`�b��|���� �$�6�_�Z�l�~�����aSSREL_IOD  �����USE_PROG %�j%�����CCRTƄ��c��_HOST !F�j! �]��T� '�y�@�R�{����_TIMEOU$��g  �`GDE�BUGƀ�k��GI�NP_FLMSK�ޟ�TR��PG��p  ���OL�C�H��yr�k�@ ����ү������C� >�P�b���������ӿ ο����(�:�c� ^�pςϫϦϸ����� �� ��;�6�H�Z߃���WORD ?	��k
 	RS�;�ZPN�q[gMAIp��SUNq���TE��ZSTsYL5r��COLXh�
��L�  ՜U�0�d�TR�ACECTL 1�
�a ��  �M�D/T Q�
��d��D � �� 5P��@��!
��"��TQ��p���PMP��IP�������	��
��U��䐾�����U�����������U�� � �  �� �7P����#�5�G�q�������Ȁ Z�l�~��������������� P�PPPP�PPPP�P��V����T�����䖆�����N���?U�F��䖾��������-?)t ����FX����U��������U�����������m��mP���������� >?Qcu��� �������� �////A/S/e/w/��/�/�/�/� I�LEpȁ]P�`�=�I�?_UP ��[Pr���q ���NQY��}d�bG_zj0�zj�&�_DEFSPD ��k{2Ђ  Т`�INPTRL ɵ���a8dU�QPE�_CONFIP�X��̈́}a��$�LIDS�����	g�LLB 1�X��P�dTB�  B4Vc}fn�Obljio��eW_ << ρ?��k�o�o�o �o �o6Nl Rd�����ZZo��=�4�a��fQ��C�����ď
eGRP� 1�;l�,�@��  �[��  � A?x�D P��DV�C2���k��E�d-�=��Q��E1���o&aY�#´��r�[�B�����������П����_a>'oY>a����K�]�G� =N�=R�b���^��� ѯ�����z��=� �xM�s�^�  Dz����_`
��ɿx�ٿ�� �#��G�2�k�VϏ� zό��ϰ������j��)Q
V7.1�0beta1_d���B(�A�?\)A�G���F��>��^����F�A���n�f�fF�A�p��AaG��q�q@�����V�� �ߵ��������p@�
�U`� #�5�G�BҢQ���� �z��v�����F�0B�ga���Ru0��e@:�� +�a��QG�@��� �� B{PB���z�BH���'�1�0��g��;Q)���x��xR�N�0n��0��R {�w���W�q�dKNOW_M ��1�c+VdSV �����U ��I[m��|�P�_b5�
cMރ��`�V�	BU����3/�CTߞ��?��@ {Q{�{Pr%n/�,�pa+MRރ��T�כּ�
��/�+̍OADB�ANFWD�+cS�Tށ1 1�Y84�Uk�V�l?_V T?f?x?�?�?�?�?�? �?�?;OO,OqOPObO �O�O�O�O�O�O_�O__572@<	!S?_`G�<}_Q_߀3g_y_�_�_574�_�_�_�_575oo1oCo57A6`oro�o�o577�o�o�o�o578*�<57MA 06��ds�WOVLD  �\{,/ȏ72PARNUM  C;���63SCH�y �u
B��P�.3b�UPD��um����U_CMP_��p���/',5ĄER_wCHK҅��,10"�Ϗ�RS� #?N�_MO ?C�_0�~�U_RES_G?0�\{
��]����� ֟���+��0�a�T� ��x���������fP����Я���P��� ��`,�K�P���_`k� �������`��ɿο�� p��υ�Xp(�G�<Lυ�V 1�F�P�	!@[l�F�T?HR_INR� �q��,5d��MASS6�� Z��MN�����MON_QUEUE �\u,6S��U�TNɀU�N
�3�J�ENDO�m�i��EXEx�iՎ�BE�w�Y�J�OPTIO�V�v�M�PROGR�AM %-�%�LІ�1�K�TASK�_I�t��OCFG� �-��!�T�D�ATA��]�~��2%�������� ���/�A�S�e�w�"������������INFO�ǡ�<ԍ�* <N`r���� ���&8J@\n������ȡ�c ��S�I�K_W���]��ENB��p�[Q&2/(G�W�2�� X,�		�=���&j/�%�!$N0���)�)���_EDIT �]��/�/P�WERFL�خ�23�RGADJ �^�*A�  55?���A5��6M���\u��?�  Bz3W��<�!����%n�?8�/W3�2Y�c7�	HD�l�ǩ��p1?� Ax�ɻt$F*%@/'B **:0B��#O�5CQM\ujBeE��AoI���?�O]M �MmOO�O�O�O/_�O �O__!_�_E_W_�_ {_�_o�_�_�_�_�_ soo/o]oSoeo�o�o �o�o�o�oK�o5 +=�as��� #��������9� K�y�o���������� ۏ�g��#�Q�G�Y� ӟ}�������ş?�� ��)��1���U�g��� �������ӯ���	� ��-�?�m�c�u�￙� ��ٿϿῦ�	p�z� �0hϡό�I��C����ϋ��&�S7PREOF �c:�0�0�
5IORITY����&�1MPDSaP��:���UT?�|C6ODUCT<���*)��6OG�_TG0A��*���HIBIT_DO�	8�TOENT �1��+ (!?AF_INE��^�~�7!tcpi�>��!ud���?!icm��>���XY\3��,��1)� =A�/��0��X�;�G���k� ������������&@8\C��*��\3�c9��?���3�>lK�7�=G/�GL�9�4��8�>A~�2,  �YЀ�����5�6)Z)�
//./�3��ENHANCOE ճ�2A�Ad(�/u%��B��J��\�11PORT�_NUM���0�x�1_CART�REP���S2SK�STA��+�SLGmS[�����3��0Unothing�/s?�?�?�<Y?��?�?�?��61TEM�P ����?8���0_a_seiban��bO��rO�O�O �O�O�O�O_�O(__ %_^_I_�_m_�_�_�_ �_�_ o�_$ooHo3o loWo�o{o�o�o�o�o �o�o2BhS �w������ �.��R�=�v�a��� ����Џ���ߏ���<�'�`�O61VER�SI������ �disable��"KSAVE ����	2670/H755J�]����!~/�����/� 	�S���:�I�|��e@��¯ԯ���J����.�9����_�� 1���|�T��������;�URGEbM B �$���WFİ ��h"��WW�崖���*WRUP_DE?LAY �>ص�R_HOT %�_Ƹ�}/e���R_NORMALD���T�<��x�SEMI�Ϯ�|��9�QSKIPd�	ܺ'u�x[�2�W�V� h�z�=�Gš߯י��� ���߹���'�M�_� q�7��������� ����7�I�[�!�� m��������������� !3EU{i����G��$RBT�IF�
<RCVT�MOU75��� DCRd���� �I�B����C4�BJ���@�/�@�I��*2T�=��]�S]¶f�� �k�����`?�a]�=ߍ��� <2�!<�"7�<L��<�`N<D��<��,�V���- /)/;/M/_/ q/�/�/�/�/�/�/�/���RDIO_TYPE  k���/�EDPROT_C_FG ��26��BHͳEE9
ѻ2�W; �8� j0�?�:��?��?�? OM�?KO��rO�ߓO ��O�O�O�O�O_�O 5_CWaOf_�-_�_}_ �_�_�_�_�_�_�_1o S_Xow_yoo�o�o�o �o�o�o�o=oBao u����� ���9>�]�� _���������ݏˏ� #�(�:���[����m� ������ٟǟ���$� C��W�E�{�i����� ï��ӯ	�/� ��G7?INT 2�Gɔ1=�AG;� ^�p��2���
Hf�0  ��Ȼ��ٯ����� B�0�f�L�vϜϊ��� ����������>�,� b�t�Zߘ߆߼ߪ��� ������:�(�^�p� V������������� �6��EFPO�S1 1�9  x�)c3�� ������*�w�����$ H��l�+� �a���2D ��+�w�K� o���./�R/� v//�/�/G/Y/�/�/ �/?�/<?�/`?�/]? �?1?�?U?�?y?OO �?�?�?\OGO�OO�O ?O�OcO�O�O�O"_�O F_�Oj_|__)_c_�_ �_�_�_o�_0o�_-o foo�o%o�oIo�o�o o�o�o,P�ot �3��i�� ��:�L���3��� ���S�܏w� ����� 6�яZ���~������ O�a������ ���D� ߟh��e���9�¯]� 毁�
����ɯ�d� O���#���G�пk�Ϳ ϡ�*�ſN��rτ� �1�k��Ϸ��ϋ�߀��8���5�n��Z�2 1�f��"�\��� �����"��F���C� |���;���_���� �����B�-�f���� %���I�������� ,��P����I� ��i��� L�p�/�S ew�/�6/�Z/ �~//{/�/O/�/s/ �/�/ ?�/�/�/?z? e?�?9?�?]?�?�?�? O�?@O�?dO�?�O#O 5OGO�O�O�O_�O*_ �ON_�OK_�__�_C_ �_g_�_�_�_�_�_Jo 5ono	o�o-o�oQo�o �o�o�o4�oX�o Q���q� ����T��x�� ��7���[�m����� �>�ُb�����!��� ��W���{����(�ß ՟�!���m���A�ʯ e���$���H���l����v߈�3 1��=�O�����+� 1�O��s��pϩ�D� ��h��ό�߰����� �o�Zߓ�.߷�R��� v�����5���Y��� }��*�<�v������� �����C���@�y�� ��8���\��������� ��?*c���"� F��|�)� M��F��� f��/�/I/� m//�/,/�/P/b/t/ �/?�/3?�/W?�/{? ?x?�?L?�?p?�?�? O�?�?�?OwObO�O 6O�OZO�O~O�O_�O =_�Oa_�O�_ _2_D_ ~_�_�_o�_'o�_Ko �_Ho�oo�o@o�odo �o�o�o�o�oG2k �*�N��� ��1��U���� N�����ӏn������ ���Q��u����4�x������4 1��� j�|���4��X�^�|� ���;���֯q����� ���B�ݯ��;��� ����[���ϣ�� >�ٿb�����!Ϫ�E� W�iϣ����(���L� ��p��mߦ�A���e� �߉��߿����l� W��+��O���s��� ���2���V���z�� '�9�s��������� ��@��=v�5 �Y�}���< '`���C� �y/�&/�J/� �	/C/�/�/�/c/�/ �/?�/?F?�/j?? �?)?�?M?_?q?�?O �?0O�?TO�?xOOuO �OIO�OmO�O�O_�O �O�O_t___�_3_�_ W_�_{_�_o�_:o�_ ^o�_�oo/oAo{o�o �o �o$�oH�oE ~�=�a�П�5 1�ퟗ� �a�L������D�͏ h�ʏ���'�K�� o�
��.�h�ɟ��� �����5�П2�k�� ��*���N�ׯr����� Я1��U��y���� 8���ӿn�����϶� ?�ڿ���8ϙτϽ� X���|�ߠ��;��� _��σ�ߧ�B�T�f� �����%���I���m� �j��>���b���� �������i�T��� (���L���p����� /��S��w$6 p�����= �:s�2�V �z���9/$/]/ ��//�/@/�/�/v/ �/�/#?�/G?�/�/? @?�?�?�?`?�?�?O �?
OCO�?gOO�O&O �OJO\OnO�O	_�O-_ �OQ_�Ou__r_�_F_��_j_�_�_o��6 1���_�_o�o yo�o�_�oqo�o�o�o 0�oT�ox�7 I[�����>� �b��_���3���W� ��{������Ï��^� I������A�ʟe�ǟ  ���$���H��l�� �+�e�Ư��ꯅ�� ��2�ͯ/�h����'� ��K�Կo�����Ϳ.� �R��v�Ϛ�5ϗ� ��k��Ϗ�߳�<��� ����5ߖ߁ߺ�U��� y�����8���\��� ����?�Q�c���� ��"���F���j��g� ��;���_������� ����fQ�%� I�m��,� P�t!3m� ���/�:/�7/ p//�///�/S/�/w/ �/�/�/6?!?Z?�/~? ?�?=?�?�?s?�?�?� O�?DO*o<d7 1�Go�?O=O�O�O�O �?_�O'_�O$_]_�O �__�_@_�_d_v_�_ �_#ooGo�_koo�o *o�o�o`o�o�o�o 1�o�o�o*�v� J�n���-�� Q��u����4�F�X� ���ޏ���;�֏_� ��\���0���T�ݟx� ���������[�F�� ���>�ǯb�į���� !���E��i���(� b�ÿ��翂�Ϧ�/� ʿ,�e� ω�$ϭ�H� ��l�~ϐ���+��O� ��s�ߗ�2ߔ���h� �ߌ���9������� 2��~��R���v��� ����5���Y���}�� ��<�N�`������� ��C��gd�8 �\��	��� cN�"�F� j�/�)/�M/�xq/WOiD8 1�tO /0/j/�/�/?/0? �/T?�/Q?�?%?�?I? �?m?�?�?�?�?�?PO ;OtOO�O3O�OWO�O �O�O_�O:_�O^_�O __W_�_�_�_w_ o �_$o�_!oZo�_~oo �o=o�oaoso�o�o  D�oh�'� �]��
��.�� ��'���s���G�Џ k�􏏏�*�ŏN�� r����1�C�U���� ۟���8�ӟ\���Y� ��-���Q�گu����� ������X�C�|���� ;�Ŀ_�������Ϲ� B�ݿf���%�_��� �����ߣ�,���)� b��φ�!ߪ�E���i� {ߍ���(��L���p� ��/����e���� ���6�������/��� {���O���s������� 2��V��z��/��$MASK 1ꊡ+����XNO  ���?MOTE  �$�G_CFG ��N��PL_RGANGJ?�%��OWER �%���SM_DRYPRG %�)��%K��TAR�T �	*UME_PRO��e/��$_EXEC_E_NB  ?��GSPD> � �(��(TDB�/�*R�M�/�(IA_OP�TION����!_AIRPUR� F*B?.�MT_� T�L2�`1g�o=�";C�?  N?�?��?�?�??1OBOT_ISOLC��>0~zENA_ME F*T/��	OB_CATEG� �O�D�uCORD_NUM� ?�;1�H755  �?�O�OY� PC_TIMEOUT�{ x� S232g�1��# L�TEACH PENDAN!Pc��pT�=JH M�aintenance Cons?�m_?"�_DNo Use�=�__��_�_oo%o�9RN�PO #R�5�6QCH_LA �̋?� 	�aso!OUD1:�ouoR� �VAIL�A5�|�1SR  /;�1��eR_I�NTVAL6��Yp> yV_DA�TA_GRP 2��� D>pP�����y �!��A�/�e�S��� w��������я��� +��O�=�_���s��� ��͟���ߟ��� K�9�o�]��������� ǯ�ۯ���5�#�Y� G�i�k�}�����׿ſ �����/�U�C�y� gϝϋ��ϯ������� �	�?�-�c�Q߇�u���߽߫����$S�AF_DO_PU�LSK�A? ��CS'CANR6�<@�SC�� �`�!X�!? �1
�2��A(�Q�U[�? ��� ���������|��#�`5�G�Y�k�HrcE�2��[��d����>	X�Hi @������?��. ��p�_ @3T01n��~�YT D��� ����"4F Xj|�������BoLe��V,/>/F$
*  =iU;�o�Tg!�EqpduE
�t��Di�@�k�Z?  � �+Jk� ��AS��/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_.a����_ �_�_oo)o;oMo_o �_���o�o�o�o�o�o��o	-2qoo0 �"�#�%�-~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N��_r��� ������̯ޯ��� o8�J�\�n������� ��ȿ3auk��� ,�>�P�b�tφϘϪ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{��������(������/�A�S� e�w�������������@��+=��
��T������"�z�	1234�5678�"h!?B!������
���f�� '9K]o��	� �����//(/ :/L/^/p/�/�/�/�/ �/�-��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO�/�/TOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_3O �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�_�o $6 HZl~���� ���� ��oD�V� h�z�������ԏ� ��
��.�@�R�d�v� 5�������П���� �*�<�N�`�r����� ����̯�����&� 8�J�\�n����������ȿڿ����"����D�V��{ύϟ���
Cz  Bp���   ���2��� }� 6��
���  	���2<�#�5�HG�Y�i���j��� ����������	��-� ?�Q�c�u����� ���������)�;�M� _�q������������� ��%7I[m��� j�k���<� ��  �������
�
�t  ���
"��`�$S�CR_GRP 1��!*P!3�0 �� ���� ��	 _m�u �k����ǒ�8��������C� ��݌*'����LR M�ate 200i�D 567890��LRMc# 	?LR2D j ��?
1234i%��x�m�� �&_ u��d�d�ӻ����)	�"?%?�7?I?[?k<��#H�u�$yd�?���?�?�?�#�����?(O�?LO�>K� �h��,Wk)�  hBB���Ɛ�O�B�D�A���O c @���E�@��@F�O ? �E�BH���_�J�F@ F�`8R@_7Od_O_�_ s_�_�_�_�_�_o� �A�AR1oo.o@oRdB�`o�_�o�o�o�o �o�o�o$H3l W�~ߥz#��w�����������A@� >ճ���@h�@U����k��' �,�;ϫ���A�@�vH΅�?�5ۀ���"��� ��*��z��M�Y�k�:�h���
 ����ß��ҟ����Y/k#DECL�VL  ������"܂A��*S�YSTEM*��V�9.10214 �s�8/21/20�20 A � �`�o�SERVE�NT_T   �$ $S_NA�ME !��P�ORT����RO�TO�� ��_SP-D��J�B�̠�TRQ   �
ɣAXISҡ�קϠ 2 �ɣD�ETAIL_ � l $DA�TETI����ER�R_COD(�IM�P_VEL�� �	:�TOQB�AN�GLESB�DIS蜠N���G��%$L�IN(� ȤREC�ҡ ,�����F�MRA�� 2w d��IDX��܋�ߠ h�$�OVER_LIM�I��栒ɣOCC�URҡ  �-�COUNTER������SFZN�_CFGҡ 4� $ENABL�(�ST"���FLA�G��DEBUF�R�[�J��Jҡ �� 
$MIN_OwVRD��$I���W�{�s���FACE��|�SAF��MI�XED�̄�d�{�R{OB��$NE��{PPôHELL ��	 5$J���BAS(�RSR�_.�  $N�UM_�B� R�1w��29�39�U49�59�69�79�98w�	�ROO��~�{CO��ONLY�p�$USE_AB����ACKEN�BA���IN۰T_�CHK��OP_S�EL_9���_PUl���M_%�OU��PNSֽ���x�9����M3�TPFWD�_KAR@���.�R�E��$OPTI{ONX�$QUE �꿠D;�Y��$CSTOPI_AL�ӆ��EX���ь�(�X�T��M1��2��M�A��STY��SO���NB��DI��T�RIFÄ�@�INIr��Mà��NRQ���END��$K�EYSWITCH�'�<����HE=�B�EATMo�PEROM_LE?�G�E<�Jn�U;�F��<�S��DO_HOM��O����EFP����Gæ�STL��C��O�M)���OV_MS��ѻ�ET_IOC#MN�Ӕ���~0���HK��
 D �-Ǳ�SU'���MP���.�PO��$F�ORC&�WARNn������OM�� �@$FU�NC� 7�U���A�R���2�3�4�~��S�O�L�Lo��!�UN�LO�%��ED�%��p�SNPXw_AS#� 0$��ADDV�X�$S�IZ(�$VAR~w�MULTIP����� Ao �� $�� ��!	&�� ��'�C;�kOFRIF��۰Sl��~	��[NF�OD?BUS_AD�&�د���CM1�DI�A]$DUMMSY1���3�4���SО� � �X�TE���8n�SGL#!TA��  &8�<#'�x� 5 $ STMT��U#PSEG��U!ByW��%$SHOW]%BANi TPO)F��9�0����SVC��Gvh� 1 $PC�ܰ� �$FBkP�(SP��A���%��VD� g�� � �A0��0�b� $1� +7� +7� +7� �+75)96)97)98*)99)9A)9B)9}  +7�+7r +7F)8�  �859��8O9	 �8i9U1v91�91�91�9U1�91�91�91�9�1�91�9���G592�B92O92\92i92�v92�92�92�92��92�92�92�92��92�93(93593�B93O93\93i93�v93�93�93�93��93�93�93�93��93�94(94594�B94O94\94i94�v94�94�94�94��94�94�94�94��94�95(95595�B95O95\95i95�v95�95�95�95��95�95�95�95��95�96(96596�B96O96\96i96�v96�96�96�96��96�96�96�96��96�97(97597�B97O97\97i97�v97c�7�97�97��97�97�97�97��97�4]�VPk�UТ ٠��.��
d V��� x? $TORu��+  D�M��RΠ��ߔQ_��R��P��G B�S��C=��F'�_U� 2����a��Lu��� �  �3ǚ
J�$0��<^��"VALU3����A�����FO�ID_YL���HI��I]?$FILE_�����$��0M�SA�ϱ hҐ�E_BLCKo�#�>!>,�D_CPU<�@<�
>����� Y# ��R  � �PW���в ��LAc!Sα������RUN_FLGŵ ��ɱ��?�̵걡�걂��Hิ���5T�2A�_LIo w �G_O��}I�P_EDI��f T2��,�4���	��7�]�  �T�BC24 �� ��̰� ��,�FT������TDC̰A��C���M�������TH�S������R��� . ERVE �������������� X -$:�LEN��G���:в�RAk��N�WI_�i�1:�פ2�דMO4��S���I���#�㡩�Ք:о�DyE�աLACE����CC�#��_M�A� ������TCV�/���T!�0�O�E�2���!s����!JJ��A�%M�䟠J��0������F�2����0����� JK��VK�!������b��J�!���JJ�;JJ�AAL��1� �1�+�
!/�5��b��N1V�b�!��!�L§�_Q!������CF�� `ҐGRO�U��?!��!N��C�S��REQUIR�EBUj6љ�7$T��2��7�p����� �� \w �f�APPR��CL�!�
$=�N0CL�Or�@	S��U	��
\��> �n�M��p�a���_MG�� C0��0	��BRK�	NOLD<�� RTMO+��
$��J+��P3��� ������O���X���%6 7 1!���� ��a��!����PATH ����f؟� ��9%�� SCAj��l1�IN9�UC�д���C0UM(Y������	!á�$*�$*:$ PAYL�OA�J2L��R'_AN��e#L��o)�k!_){!�R_F2�LSHR	Ԩ!LO�p$��'#�'#ACRL_y��� �W$rY�H��!�$H��2FLEX3�:��J�� P�ϐ��� ߞ�319�  :F�X��Щ7��4[�Z���d�v߈�F1�1E"G�ߩ߻�������RBE����1� C�U�g�y��)XFT�� ����6@XX�����1��T�W'QX�0Q�� �D}H���U�H���� 0�4�=�+�O�X�j�|�p����40��! ���`����������AT;F���EL�@�s���J�� ��JE� C3TR�6ATNƑ	v���HAND_VB�!�31��t" $��PF2�����S�W�����~#� $$M� �	����x��|�@�u�vA@Ơ\ �š��A����
A�A���TU��
D�D�P�G����ST����	��N�DY˰. � �t�} ;П'�1�'�!@^'��}T�0�P�P( 1:CLU^g�2�t$ �p�4� �cA��b��ASYIM�#����#���!�_��(�$ ����x/-/?/Q/c#Jj,|*�����)HD_VIds٨b�V_UNK�ؠ�� c�!J���E���,� �%(�L��-���)�/?���S$4,3l��3HRt�i�%zrͱLF0@�DI� ��O��  �ͱ�c&) 0`�I�A�#��<@'�'�?@p����Aϰ ' � -�qME�At`B�4��)�T�PT��`�j���dE0a�o���~�T���� $DUMMY1:�$PS_9@RF��0l$��� FLA��YP�S��r�$GLB_T�p ���j�N1�0x@:qF��( X ��tST��A��SBR�M�21_V��T$S/V_ER� O��@ӦX�CL�@�A�@Ol�ɰGL�EW���) 4��t�$Y
qbZqbW����!�s�AC�" ��U.��* �PN�Ѕ��$GIJp}$��� �ЃӼФ�+� L����S�}$FzS�E��NEAR�@�N@CF-�@TAN9C@BlJOG�0� ,��$JOgINT�Q�PC_���MSET��-  "��E�A�`S�b��|�a��.� Bp�U�A?���LOC�K_FO� �q�B�GLV=sGL��T?EST_XM3 ��'EMPi�����Ҏ��$U�0���P2*���!�+��p��!�)B�CE����B�_ $KAR�AM�TPDRA��_�V��VEC�0p�Z�IU�!�,&�HE��TO�OLC��VDRENw�IS3�5��6CN6@ACH|���-��QO�rô�30a���SI#  @$�RAIL_BOX�E�Qe�ROBO���?�e�HOWW�AR1����ROLM��7�a��H�a���*@vO_F�`!}e�HTML5�j�ƳGJ CHw�/b���Rz�OB�20b��0k�o ��v��OU~�1 d����))�r�a��$PIP��N�P�������H@!� �0COR�DED���� *�XIT� ��)ɰ�`O)� 2 D ��OBE�s��P?��p��?S�qSYS?�ADRqɰj�TC}H�p 3 ,�PSENҲO1A��_�Ա��a'�ACɰV�WVAE�4 �� e����PRE�V_RTR�$E�DIT�VSHW�R�a,� �B���٠DT��1'$ a$HEADd���A �t��KE�Ѩ�C�PSPDX&JMP�\L���R�@�Q5GD1�I��Sr�C^pNE��qTwT�ICKC�MM1�s�#HN"�6 �@I�!�e`!_GP8�&��P0STY���LO�hr�"�"�0_7 t 
�G�S%$���=,�S`!$��PY����r��P��&SQUY�x�5��ءTERCn��N��TS�d8 ��8��g�P�g%Q��b)�Oo�b�D@IZ��4������PR%���B�!� PU�aE_�DO2�XSz�KN�AXI<@[&�UR�`�Cr � jd�q�`_��|ET}BQP��Xҕ;0Fҗ�<0A߁Ց��9���)��ƲSRqt9l�0�y�R�z�E �v
Y�r�E�w�C��C �>U3�>UC�>US�PU@j]��PU�\��nYC�_|]C�]L�^�p�����SSC�� : �he�DS� `��S�P�jeATA��r�A� �"��ADDR�ES��B�SHIyF�c�_2CHp�fIмa�TU��I�q ;b�COUSTO�D��V��I�<���~aC��
��
�V�-AG�'= \*���;0|�1�0IrC��2�Bz��^�Iq�TXSCWREEA>ٰW1TINA{��Мt���}!~A~b��? T �![�B|Z�7��vJAp{JB�t�RRO��G�{R �q8���UE��$@ ������S�|�|RSM� @GU`.�0�S�ͰS_�Ӏs��c�v����~ACx��O��t 2?�pUE��A�kҶ�@WGMT_�L9�YA�G�Ol�'0BBL_r��W��G�B �;0j�O���LE�b�*� �b)�RIGH�3�BRDmԤaCKGR��[�T/Z�W�WIDTH�� 7¨������2�Ij E	Y~`F�C�z 6 2z��	ABACK1h��Εq�M�FOn�LAB(Q?(M�yI����$UR��S৐S�H	� 'D 8��G�_@!�b1�T�R�����C��������O�aG�E� $x�T�U?��R��B�LUM�aF�`ER�V��Ч�P1ஔFK��@GE��@L5I LPѥ�BE�0/a)�?a��Oa������5��6��7��8 ޢ�2b�@1�]t������S�0E��U{SR��G <*�bS�U���c��FO�`.��PRI�Am��m��аTRIP��m_�UNDO�H���`0�BE)AE��8�{@u0 I,���.AG H0T[ aL�a'�OSr�<�R�@�Û�ӁJ�ߤӫސc��$ˁ�U١ӁK�l�~ό�٢�%�OF�F����L(���OD��"�Je����Ke�GUvPѬB�a)׻�SUB�"tТ�RTe��DM�"F�g ��3OR��o�RAUD�@p�T�٢U�_�·$N |�@�OW�N��$SRC����^0D�����BM�PFI4a}@ESPA�2�p����.!���� ��
 ӁO `&��WO$P��1�07COP��$r@��_�м�i��p�WA�C��M�#�L��p'0�5�a P�r?SHADOW^@��~��_UNSCA~�8�㓔��DGD��W�EGACc�w��VC P)�ӁQ�c ��@l3$��ER�p,��1����C�� ,�DRIV�6��A_V� O�� 6 D~|�MY_UBY{� 4�B6c�l5��0�p.!1��1���P_��4���L#KBM&�$n� DEY�EX �,'�t�MUv X&��h�US]�h@˰_R@�q�����`���G�P�PACIN�!i0RG��Xn��n��n��i�REF��ac��Bq�n�R �`
[�Gt�Pr� ���	RS��S��x�����O�	h�:ARE+SMWf _Ag�@ @O���aA�`'�BEEl�U.0H��A�V�HK32Tu�?`���A$�ppEA� �zL�3�'��MR�CVӁU �ʠO*?0M3�C�s	�����REF���� ����C� ���!@�!�1%�f_��|g(�xPSi�����1{1Z��ЄV �@2�����0�����0�OU�'��&4� SQ�a2��$�p_p@��S}ca�!lD��`UL�pT(�3COG�H�U 0NT#�P41�O5`�[6��[30L��5��5�`��7���VIA�_L�]`W ��@HyD�`Ɛ$JOg�����$Z_USPL̰ �ZEPW�5p�139���_LIM�$EP1I�4��1 �1�q�a���`
�0&�>6�X� 0}c�Az@` }cCACH��LO!lD�A �I���|���C@MI�cF�A�ETVP�F�+$H�O3���p@COM	MJ�O�O=��G�'��`d3��͡�$ �VP�<��6R_SIZ��@T�ZR ;X�1<W��n�M]P`ZFAI�0Gl��@AD�Yi�MR1E�$�REWGPU� ���s�ASYNBU=Fs�VRTD�U�TlEQn�OL�`D_���
eW��PC�`TU� �@QD�UECCU�VEM� �ERb�GVIRC�Qe�S|N��Q_DELA�����簶�AG�YR�XYZ��}�W@��h!�d��o`T�IM�af�b���E_GRABB`�Y+�� %�ЄY��ڒL�AS���PA_GE�WEZ>���sbc_uT@�#���)����I�tX��fb�BG/�V���p�PKq �fXA�'GIOpN�)R�Kq�@$�Q:�[���AS�P}F�N��LEXPv\���ӳ��z�Q��I  �S��E���E���mE֐��b����]���+��DY�����*�ORDı�{�°@��"��^ $0TIT��ɰ������VsSFv���_  ���$�[1 UR��PS�M�`����AD�J΀�0ZD�a3 D��AAL�0�P<Π
BPERI<@���MSG_Qc$@FQdU[���eBa�b��`�0�@���@�W�XS�h�c��� uK�CH)�HOL��]��XVR�d7r�+�T_OVR2�_�ZABC\�e��6��C�
MAc�z�V�S@ f � �$_��|�CTIVz��AIO���FfY�IT
�mDV	�#
mX@��{Q��MàPS�!�� �S����A� ���ALST`Y��A�00��_S���$qc�DCSCH��g Lg�#�w���@ �GÀ@� EPGN�A�C���A"�_F#UN��@��Z&�촙h���$L����  �ZMPCEF\�i���
���f��LN ��
@����`]�j $x�Az��CMCM` ECr�C\����P^�? $J��D+Q!�2�+ǚ07Ś0`Ǩ��0�c�UX�a��UXE&���a&� z�<�z����Ɍ����FTF<1!�������k D��������Y@Dp l� 8cR�PU��?$HEIGHY�#?(0ؖ����>�$m � �S��$B0A���L�SH�IFvS��RV@F�����+�C�0�\� -4�D��ְ^s�� UYD���CE��V}!}m��SPHERh� n ,00�F�fX��r���FA;1��c���u�{�S�HOT��_��@S�MIPOWERFL y��c�k� ��WFD�O`� ��G@� 1� ������� L!��_EI�P���c��j!�AFz0E_�$���!'FT��S��w�3!�x����f���7!R'`MA@����������p��������[!OPC3UA\�
J�!TPz0p���yd��!
PM�&�XY��e�?Ⱥ	�f.�!�RDM�V��g|z�!R90�2	�h�#/!
���@�X�i/o/!ReL�PCp/�)8^/>�/!ROS���,��4�/?!
CEF� MT�@?�k�/S?!	2C{�q?��lB?�?!2WA'SRC��m�?�?;!2USB�?��n�?7O!STM��QO�o&O�O���OКtO�M��I
�KL� ?%�� (%�SVCPRG1��OZU2__P3�@_E_P4h_m_P5��_�_P6�_�_P7��_�_P8ooP90o5kT�]oQ
_ �oQ2_�oQZ_�oQ �_�oQ�_%Q�_M Q�_uQ"o�QJo �/Qso�/Q�o�/Q �o=�/Q�oe�/Q�� /Q;��/Qcݏ/Q� �/Q�-�/Q�U�WQ ��O�BG`�O P��� 'Q����1��U�@� y�d�������ӯ���� ���?�*�Q�u�`� ���������̿�� �;�&�_�Jσ�nϧ� �Ϲ��������%�� I�4�m��jߣߎ��� ���������!�E�0��i��J_DEV ����MC:�t��GRP 2���� �@bx 	�� 
 ,�� q��﬒�����9� � 2�o�V���z������� ����#
G.k }��X���� �1U<y` r�����	/� -/�"/c//�/n/�/ �/�/�/�/??�/;? "?_?q?X?�?|?�?�? �?�?F/O%OOIO0O mOTOfO�O�O�O�O�O �O�O!__E_W_>_{_ b_�_�_O�_�_�_o �_/ooSoeoLo�opo �o�o�o�o�o�o+ =$a�_V�N� ������9�K� 2�o�V�������ɏ�� �ԏ�#�zG�Y�@� }�d�������ן���� ��1��U�<�y��� r�����ӯ�<�	��� -�?�&�c�J������� �����ȿڿ���;� "�_�q�Xϕ�쯊��� �������%��I�0� m��fߣߊ������߀����!���W��d �^�	E��y��`��������	�%�	�<.������G��� G�W�e�O���s����� ����� C���- Q?acu���� ��)M; ]������� /�%//I/�p/� 9/�/5/�/�/�/�/�/ !?c/H?�/?{?i?�? �?�?�?�?�?;? O_? �?SOAOwOeO�O�O�O �OO�O7O�O+__O_ =_s_a_�_�O�_�_�_ �_�_�_'ooKo9ooo �_�o�__o�o�o�o�o �o#G�on�o7 �������� aF���y�g����� ����я'�M��]��� Q�?�u�c��������� �#������'�M�;� q�_���ן������� ݯ��#�I�7�m��� ��ӯ]�ǿ���ٿ� ���Eχ�lϫ�5ϟ� ���ϱ������M�2� D������eߛ߉߿� ����%�
�I���=�+� M�O�a�������� !����9�'�I�K� ]������������� ��5#E����� ��k����� 1sX�!�� ����	/K0/o �c/Q/�/u/�/�/�/ �/#/?G/�/;?)?_? M?�?q?�?�?�/�?? �?OO7O%O[OIOO �?�O�OoO�OkO�O_ �O3_!_W_�O~_�OG_ �_�_�_�_�_o�_/o q_Vo�_o�owo�o�o �o�o�oIo.mo�o aO�s��� 5�E�9�'�]�K� ��o����̏����� ���5�#�Y�G�}��� ���m�ןş���� 1��U���|���E��� ��ӯ������-�o� T������u�����Ͽ ���5��,���߿ Mσ�qϧϕ������ 1ϻ�%��5�7�I�� mߣ�����	ߓ����� !��1�3�E�{�ߢ� ��k����������� -����z���S����� ��������[�@� 	s����� �3W�K9o ]����/ �#//G/5/k/Y/{/ �/��//�/�/�/? ?C?1?g?�/�?�?W? y?S?�?�?�?O	O?O �?fO�?/O�O�O�O�O �O�O�O_YO>_}O_ q___�_�_�_�_�_�_ 1_oU_�_Io7omo[o �oo�o�_o�o-o�o !E3iW��o ��o}�y��� A�/�e�����U��� ���я���=�� d���-���������ߟ ͟��W�<�{��o� ]���������ۯ�� �˯�ǯ5�k�Y��� }�����ڿ������ ��1�g�Uϋ�Ϳ�� �{�����	����� -�cߥϊ���S߽߫� ��������kߑ�b� ��;��������� �C�(�g���[���k� ���������� ?� ��3!WEg�{ ������/ SAc���� y��/�+//O/ �v/�/?/a/;/�/�/ �/?�/'?i/N?�/? �?o?�?�?�?�?�?�? A?&Oe?�?YOGO}OkO �O�O�O�OO�O=O�O 1__U_C_y_g_�_�O _�__�_	o�_-oo Qo?ouo�_�o�_eo�o ao�o�o)M�o t�o=����� ��%�gL���� m�����Ǐ��׏��?� $�c��W�E�{�i��� ��ß������՟�� �S�A�w�e���ݟ¯ ���������O� =�s�����ٯc�Ϳ�� �߿���Kύ�r� ��;ϥϓ��Ϸ����� ��S�y�J߉�#�}�k� �ߏ��߳���+��O� ��C���S�y�g��� �����'���	�?� -�O�u�c��������� ������;)K q�����a��� �7y^p' I#�����/ Q6/u�i/W/y/{/ �/�/�/�/)/?M/�/ A?/?e?S?u?w?�?�? ?�?%?�?OO=O+O aOOOqO�?�?�O�?�O �O�O__9_'_]_�O �_�OM_�_I_�_�_�_ o�_5ow_\o�_%o�o }o�o�o�o�o�oOo 4so�ogU�y� ���'�K�?� -�c�Q���u����ҏ 䏛������;�)�_� M���ŏ���s�ݟ˟ ���7�%�[����� ��K�����ٯǯ�� ��3�u�Z���#���{� ����տÿ�;�a�2� q��e�Sω�wϭϛ� �����7���+߽�;� a�O߅�sߩ������ �����'��7�]�K� ���ߨ���q������� ��#��3�Y������ I������������� a�FX1y� ����9]g��$SERV_M�AIL  g�]�COUTPU}TRh }@GRV 2�;  ` (�-<�GSAVEsa�TOP10 2>� d c/ +/=/O/a/s/�/�/�/ �/�/�/�/??'?9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O0�O_��YP�D�FZN_CFG ;�`$���MQGRP 2�WW� ,B �  A�PgD;�� B�P�  B�4#RB21��HELLPR	����nW ok%RSRoo"o [oFoojo�o�o�o�o �o�o�o!E0i�{�~�  ��]r����r� �h ��r�q�x�r2�h d�|�}8��VHKw 1
�[ � r�|�v���ɏď֏� ���0�Y�T�f�x�࡟�������\OMM� �_��RFT?OV_ENBR���P�OW_REG�_UI0�EIMI_OFWDL������Ue�WAIT-� 1�oR��mQ����wTIMQ���į�VAQ��e�_UNcIT,����LCJ�WTRYQ��G�MON_ALIA�S ?e���he�������úm� ���
��ǿ@�R�d� vψ�3ϬϾ������� ���*�<�N�`�߄� �ߨߺ�e������� &���J�\�n���=� �����������"�4� F�X�j���������� o�����0��T fx��G��� ��,>Pb s����y�/ /(/:/�^/p/�/�/ �/Q/�/�/�/ ??�/ 6?H?Z?l??�?�?�? �?�?�?�?O O2ODO �?hOzO�O�O�O[O�O �O�O
_�O_@_R_d_ v_!_�_�_�_�_�_�_ oo*o<oNo�_ro�o �o�o�oeo�o�o �o8J\n�+� ������"�4� F�X��|�������]� Ï�����ɏB�T� f�x���5�����ҟ� �����,�>�P�b�� ��������g���� �(�ӯL�^�p������>��$SMON_�DEFPROG �&������ &*S?YSTEM*��߷�p��?��R�ECALL ?}��� ( �}:�copy frs�:orderfi�l.dat vi�rt:\tmpb�ack\=>16�9.254.E�1�20:17084�߿e�wφ�}1�m?db:*.*/�Aσ4 L�����ߔ�5x�:\��$е��°��a�s߅�}6�a�"�4�K�Q����߇�
�xyzrate 11 �߷���Z�l�4~��!�24:�P� ��N���������+� ����`�r�����2��� M������(��K� \n���$6��� ���#���G�Xj |����<����� �CT/f/x/���./�S/�/�/��� �/�/�/[?m??� ��E4964� ;?M?�?�?O�9 ,�?�1SOeOwO�0�5O�:KO�O�O _�4/-?�>�O`_r_ �_(�/3_�7P_�_�_ o?�_�_�__oqo�o<�?�;6640�>Ko��o�o �tpdisc 0�o�a�o��o[m�tpconn 93E ���OO�O�nS� e�w��O�O7��hK�܏ � �_&o8o�cϏ`� r����_(�:�L�Q�� ����﫟��ϟ`�r� ���o>���M�ޯ�� �����ɯZ�l�~��� ��5�G�ؿ����!� ��ſV�h�zύ���1� C������������� �d�v߉���6߿�Q� ���߇��,�����`� r�(�:������� ��'߰���\�n��� �ߥ�@�����������$SNPX_A�SG 2����%� � ��%�M � ?�PARAoM %/� �	;PrP��& � OFT_KB_?CFG  +�OPIN_SI�M  %���( RVN�ORDY_DO � ��:QS�TP_DSB���~SR �%	 � & �LABWELD_�2����T�OP_ON_ER�RG�PTN �% ��A	"RING_P�RM�YVCNT�_GP 2��2 x 	zy/�g/��/�/�/VDN ROP 1u	� �! %�/�/?#?5?G?n? k?}?�?�?�?�?�?�? �?O4O1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_o�o�o�o�o�o �o�o�o%LI [m����� ���!�3�E�W�i� {�������؏Տ��� ��/�A�S�e�w��� ������џ����� +�=�d�a�s������� ��ͯ߯��*�'�9� K�]�o���������ɿ �����#�5�G�Y� k�}Ϗ϶ϳ������� ����1�C�U�|�y���ߝ߯������"PRG_COUNT�s�"��ENB4/���M$��1�_UP�D 1�T  
���{����� ���������/�X� S�e�w����������� ����0+=Ox s������ 'PK]o� �������(/ #/5/G/p/k/}/�/�/ �/�/�/ ?�/??H? C?U?g?�?�?�?�?�? �?�?�? OO-O?OhO cOuO�O�O�O�O�O�O �O__@_;_M___�_ �_�_�_�_�_�_�_o�o%o��_INFO� 1i�O�q`	 Ho�owo��o�i?�̬@d��7=��?q{*�o B�;c�7���o�g>C�P ?�2 A6�~��b�n >���{ �'���Dd�8C���6���X ��b@p�d�����XD̿7�3���W����3���YSDE�BUG	�j��?`d�R�zpSP_PAS�S	�B?�{LO�G ffs� � ?`xEo  ��aq`  UD�1:\�tLn�r_M�PC�}i�:�L�i���o>bi��SAV �y�a�q�r;e� �SV�TE�M_TIME 1u�wt� 0O�aWK��L�l� ʇ�MEMBK  i�N��p�N�`�p��X|O�� @p�;cВ���ǜ��d�����q �k@�/�A�S�e���}��������ůׯ� � ��!�3�E�W�i�{�������e��ӿ��� 	��-�?�Q�c�uχ� �ϫϽ���������)�̅SK%�*��9��i�{ߍ߁�4?`X�,�2����A��p �� ֒"��� ���$�T�f�ʟl���  �����;c����������߀+�P�b�t�����?`$������ ����,>Pb t��������(:.�T1SVGUNSPD�u� '�u�]2M�ODE_LIM !,�恐rY2f���}XASK_?OPTION�p-���q�_DI�pENB  ���u��BC2_GRP 2LՌs�$/����C�9#QBCCFOG +����p*`�/�o�/�/ �/�/�/ ??D?/?h? S?�?w?�?�?�?�?�? 
O�?.OO>OdOOO�O sO�O�O�O�O�O_�� �L _�OS_e_�OB_�_ �_�_�_�_q�o/��P o1ooUoCoyogo�o �o�o�o�o�o�o	 ?-cQs��� �������)� _�E�0Ps�������Ǐ E��ُ��!��E�W� i�7���{�����՟ß ����/��S�A�w� e�������ѯ����� ��=�+�M�O�a��� ����q�ӿ���'� ��K�9�[ρ�oϥϷ� �ϗ��������5�#� E�G�Yߏ�}߳ߡ��� �������1��U�C� y�g��������� ���ѿ3�E�c�u��� ����������� )��M;q_�� �����7 %[Ik��� ����//!/W/ E/{/1��/�/�/�/�/ e/?�/?A?/?e?w? �?W?�?�?�?�?�?�? OOOOO=OsOaO�O �O�O�O�O�O�O__ 9_'_]_K_m_o_�_�_ �_�_�/�_o#o5oGo �_koYo{o�o�o�o�o �o�o�o1UC egy����� ��	�+�Q�?�u�c� ��������͏Ϗ�� �;��_S�e������� %�˟��۟��%�7� I��m�[�������� ůǯٯ���3�!�W� E�{�i�������տÿ �����-�/�A�w� eϛ�Q���������� ��+��;�a�O߅�o�����$TBCSG_GRP 2o���  ��� 
 ?�  ���������(� �$�^�H���Ү����d@ ����?��	 HBL������B$  �C�����	�����C�z	�Q�AД�33�3?&ff?�����A����a� ����ͷ�|���DH����@�q��t� ����D"w��� ��d/
��r��� �u������:Ic	V�3.00��	lwr2dI	*�0}�ҔS �� ���  ��/+��J2����fG/$%CFG [!o��� ��K*�u"�x,�,��/�/�*x��/ �/�/?	?B?-?f?Q? �?u?�?�?�?�?�?O �?,OO<ObOMO�OqO �O�O�O�O�O�O�O(_ _L_7_p_�_�����_ �_�_[_�_�_�_oo >o)oboMo�o�o�o�o wo�o�o�o:�� ��_k�oq��� ����%��5�[� I��m�����Ǐ��׏ ُ�!��E�3�i�W� ��{���ß���՟� ���5�G��g���w� ����ѯ������+� =�O��_�a�s����� Ϳ߿�Ͻ�'��K� 9�[�]�oϥϓ��Ϸ� �������!�G�5�k� Yߏ�}߳ߡ������� ���1��U�C�y�g� ���Y��������� 	�+�-�?�u�c����� ����������; )Kq��O�� ���7%G I[����� ��/3/!/W/E/{/ i/�/�/�/�/�/�/�/ ??A?S?��k?}?;? 9?�?�?�?�?O�?O O+OaOsO�OCO�O�O �O�O�O__'_9_�O ]_K_�_o_�_�_�_�_ �_�_�_#oo3o5oGo }oko�o�o�o�o�o�o �oC1gU� y����_?�� !��Q�?�a���u��� ��Ϗ�����)�� M�;�q�_�������˟ ������%��I�7� m�[�}�����ǯ��� ٯ����!�3�i�W� ��{�����տÿ�� ��/��S�A�wω�3� �ϳ�9�o������� =�+�M�s�aߗߩ߻� yߋ�������9�K� ]�o�)������ �������5�#�Y�G� i���}����������� ��UCyg ������� ����EW/u� ����/�)/;/ M/_//�/q/�/�/�/ �/�/??�/7?%?[? I??m?�?�?�?�?�? �?�?!OOEO3OUO{O iO�O�O�O�O�O�O�O �O_A_/_e_S_�_w_ �_�_i�_�_�_�_+o oOo=o_oaoso�o�o �o�o�o�o'K89oY~  �p�s� �v��r�$�TBJOP_GR�P 2"au��  ?�ҙv	�r�s$�|��ip�@�� 0�u � � � � ߈ ��t �@�p�r	 �B�L  I�Cр D�w�qe�>�n�j�~|�<�B$?�����@��?�33C�S���a����ǇI�[�}����;��2������@_��?��z;����V�A�g��〝a ���6��p>̧�|����;��pA:��?�ff@&ff�?�ff��ޟa� ���u�󄦁��,�:7v,���?L�����ʐDH�^�d�v�@G�33����>ʐx������8��퉡�q=�2�D"������������=�9�K�9��ݯ﯐����� ��חɿ����� ��� ��?�Y�C�Q�ϰϋ� E����������@ߙs�C��v2���	�V3.0�	l7r2d�t*���t��q�ߤ� E8�� EJ� E\� En@ E�p�E�� E�� �E�� E�� �E�h E�H �E�0 E� �Eϻ��� E����� E�x E�X F����D�  D�` �E��P E���$��0��;��G���R��^p Ek���u����І���(��� E��Н��УX 9�IR$]�)�q������
���v��9�՟����tESTPARS�r��x�p�sHR��A�BLE 1%�yJs��t��� `��������w�q*��	��
����.�*�q������t�N�RDI��q-�@?�Q�c�u�����O���	%7I[�S���s ��.@R dv������ �//*/</N/`/r/ �}� ��r,��)�� ��~�������������"NUM  Vau�q%��p� s�t��_CFGG &�;/3=�@�p�IMEBF_TT���*5�s��6VER�r��!�6�3R 1='� 8�ߙr��p7A dp�/   O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_�_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[� ������� �!�3���A_|1�6�@�5��MI_CWHAN�7 �5 ���DBGLVڀ�5��5�ᡀETHER_AD ?������G�E�����ޡ�ROUT�0!ƀ
!S�q�D�SN�MASK��3��255.��wӭ����џw���OOLOF/S_DI��k�Ӊ�ORQCTRL C(Kg��O�T>� s���������ͯ߯� ��'�9�K�]�o��������=�ƿ�����PE_DETAIǈ��PGL_CON?FIG .�9�1���/cell�/$CID$/grp1�d�vψϚ���b�:�������� �1���U�g�yߋߝ� ��>�������	��-� ����c�u����� L�������)�;��� _�q���������H�Z����%7I�.} �������G1ۿ����6HZ l~������� �/�2/D/V/h/z/ �/�/-/�/�/�/�/
? ?�/@?R?d?v?�?�? )?�?�?�?�?OO*O �?NO`OrO�O�O�O7O �O�O�O__&_�OJ_ \_n_�_�_�_�_E_�_ �_�_o"o4o�_Xojo |o�o�o�oAo�o�o�o�0B=���User Vie�w R�}}1234567890s ������t^�2����Yy2fy�o7� I�[�m������`r3�ߏ���'�9���Z��4Ώ������@ɟ۟�L���5�� G�Y�k�}����� �¯�66�����1�C�U���v��7꯯����ӿ���	�h�*��8 ��c�uχϙϫϽ������� l?CameradzZπ#�5�G�Y�k�}�[E ߧ߹���q����	�0�-�?�5�  ��� ߏ���������� ��1�|�U�g�y������������͉F��� 1CU��y� �������	 �������gy�� ��h��	/T-/ ?/Q/c/u/�/.��[�  /�/�/�/??/?� S?e?w?�/�?�?�?�? �?�?�/��驊??OQO cOuO�O�O@?�O�O�O ,O__)_;_M___O �����O�_�_�_�_�_ o�O)o;oMo�_qo�o �o�o�o�or_��Q�bo );M_qo� ������%�7��o�g9�x����� ����ҏy���� +�P�b�t�������9�	��00����	�� -�?��c�u���.��� ��ϯ�������� ۩�^�p��������� _�ܿ� �K�$�6�H� Z�l�~�%���r���� ���� ��$�˿H�Z� l߷ϐߢߴ������� ��˕����6�H�Z�l� ~��7ߴ�����#��� � �2�D�V����J ���������������  2D��hz�� ��i��+Y  2DVh��� ����
//./� �"K�z/�/�/�/�/ �/{�/
??g/@?R?�d?v?�?�?A-  E)�?�?�?�?O#O�5OGOYOkO}O�K   �?�?�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q�����p����L  
A �(  �0( 	 �G�5�k�Y� ��}�����Ïŏ׏����1��U���J ��/������1?� ����*�<�C#��f� x���џ����ү��� �O�,�>�P���t��� ������ο���� ]�:�L�^�pςϔ�ۿ �������5��$�6� H�Z�l߳ϐߢߴ��� ������� �2�y�V� h�z��ߞ�������� ��?�Q�.�@�R���v� ������������� _�<N`r�� �����%& 8J\����� ����/"/4/{ X/j/|/��/�/�/�/ �/�/A/?0?B?�/f? x?�?�?�?�???�? OOa?>OPObOtO�O �O�?�O�O�O'O__ (_:_L_^_�O�_�_�_ �O�_�_�_ oo$ok_K�@ FbSoeowo�FcMg1���+f�rh:\tpgl�\robots\�lrm200id~�`_mate_�b.xml3o�o�o %7I[moV�������� ��,�>�P�b�t�� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l���}�����Ư د���� �2�D�V� h��y�����¿Կ� ��
��.�@�R�d�{� uϚϬϾ�������� �*�<�N�`�w�qߖ� �ߺ���������&�8�J�\�n�h�Q� Mo�`<< �` ?�n��n� ���������/��G� e�K�]���������� ������3aoV��$TPGL_�OUTPUT �1yQyQ �������� 0BTfx� ������//�,/>/P/����f 2�345678901u/�/�/�/�/�/�# oRr/�/?"?4?F?X? �/\?�?�?�?�?�?n:}�?OO,O>OPO�? �?�O�O�O�O�O�OxO �O_(_:_L_^_�Ol_ �_�_�_�_�_t_�_o $o6oHoZoloozo�o �o�o�o�o�o�o 2 DVh ��� �����.�@�R� d�v��������Џ� 􏌏��*�<�N�`�r� �������̟ޟ�� ���8�J�\�n����q}�ᶯȯگ�����!�@��E�W���? ( 	 Z/�� z�����Կ¿���� 
��R�@�v�dϚψ� �Ϭ���������<� *�`�N�p�r߄ߺߨ���h&�������*� �L�^�8���b*�� ����q��������C� U���Y���%�w����� ����	g���?��+ u�a���� �);Gq� ���S���� %/7/�[/m//Y/�/ }/�/�/�/I/�/!?�/ ?W?i?C?�?�?�/�? �?�?�?OO�?%OSO �?;O�O�O5O�O�O�O �O_eOwO=_O_�O[_ �___q_�_�_+_�_o �_�_9oKo%ooo�o�_ io�oQo�o�o�o�o# 5�ok}�� ���GY�1�� 9�g�A�S������ӏ ��я����Q�c����)WGL1.�XML!����$T�POFF_LIM� ��+�������N_SV�� � (���P_M�ON 2���+�+�2��ST�RTCHK 3���������VTCOMPAT՘_�Ė�VWVAR 4r����ٔ 6�� �������_�DEFPROG �%$�%MA�IN ELD_1�����_DISPL�AY��$�ʢINST_MSK  �� �INUSsERU��LCK^��%�QUICKMEyN���SCRE�����`�tpsc�^�������Ұ�_ֹSTS���RA�CE_CFG U5������	���
?��HNL C26٪��A��� �� uχϙϫϽ����������ITEM 2�7a� �%$1�23456789y0H�Z�  =<R�xxߊߒ�  !���۬�\��ߣ�F�� j�*�<��R����ߟ� �ߺ������v�f�x� ����(���~����� ���>�P�b�����2 Xj��v��� �L�*�� ��� ��6� Z�5/�P/�`/�/ �/��/ /2/D/�/h/ ?:?L?�/p?�/�/�/ |?�?.?�? Od?O�? �?cO�?~O�?�O�OO �O<ONO_rO2_�OB_ h_�O�O�O__&_�_ J_�_o.o�_Ro�_�_ �_To�_�o�o�oFo�o jo|o�o`�o�� �o�0�T�x 8�J��`��$���� ȏ,�؏���t���� ����6�������ğ(� �L�^�p������f� x�ܟ�� ��ۯ6��� Z��,���B���Ư����S'�8-ϔ��g  Ҕ� 9���
 �����B�úUD1:\�O�����R_GR�P 195�� 	 @렚Ϭˀ���Ϻ������ޠ $�;�I��O�s�^ߗ���?�  ���ۮ� �������,��<�>� P��t�����������(�	b�<�N�~��SCB 2:�� �ߚ������������*��UT�ORIAL ;�6�u��V_CONFIG <���4��2���OUT?PUT =��� ���$6H Zl~����� ���$/6/H/Z/ l/~/�/�/�/�/�/�/ �// ?2?D?V?h?z? �?�?�?�?�?�?�?	? O.O@OROdOvO�O�O �O�O�O�O�O_O*_ <_N_`_r_�_�_�_�_ �_�_�_o_&o8oJo \ono�o�o�o�o�o�o �o�oo"4FXj |������� �0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ����P� b�t���������ο� ���(��L�^�p� �ϔϦϸ������� � �$�5�H�Z�l�~ߐ� �ߴ���������� � 2�C�V�h�z���� ��������
��.�?� R�d�v����������� ����*;�N` r������� &8I\n� �������/ "/4/EX/j/|/�/�/ �/�/�/�/�/??0? A/T?f?x?�?�?�?�? �?�?�?OO,O>OO? bOtO�O�O�O�O�O�O��O__(_:_����Y_k_UQD_�_ 9��_�_�_�_oo&o 8oJo\ono�o�oEO�o �o�o�o�o"4F Xj|���o�� ����0�B�T�f� x��������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϯ������� ��
��.�@�R�d�v� �ߚ߽߬�������� �*�<�N�`�r��� �����������&� 8�J�\�n�����������$TX_SCR�EEN 1>mU�UP�}������	-?Q ���V������� �bt!3EWi {������ //�A/�e/w/�/ �/�/�/6/H/�/?? +?=?O?�/s?�/�?�? �?�?�?�?h?O�?9O KO]OoO�O�O
OO�O �O�O�O_#_�OG_�O k_}_�_�_�_�_<_�_��$UALRM_�MSG ?����� �_��o-o^o Qo�ouo�o�o�o�o�o� �o$H�USEoV  
mzv��RECFG @v����  ���@�  A�q  w Bȶ�
 I ��������%�7��I�[�m�������qG�RP 2A�{ 0��	 ���P�I_BBL_NO�TE B�zT?��l�������p��DEFP�RO`%
k (%<c���Q���u��� ��ҟ������,���P�;�t��FKEYDATA 1C���Ӏp �w���֏ٯ�¯�!���,�(-�T���(PO?INT  ]\�^��WELD_ST�������P��߿��E�ND��TOU�CHUP��  �ORE INFO 8�;�xϊ�qϮϕ��� �������,�>�%�b��I߆ߘ� ���/frh/gui�/whiteho?me.png���߰��������point��S�e�w����*���arc_strA�E��������'����weldB�]�o�������4���enK������(��touchup��ew���:����wrgA�� �/��8\n ����E��� /"/4/�X/j/|/�/ �/�/A/�/�/�/?? 0?B?�/f?x?�?�?�? �?O?�?�?OO,O>O �?POtO�O�O�O�O�O ���O�O_ _2_D_V_ ]Oz_�_�_�_�_�_c_ �_
oo.o@oRo�_do �o�o�o�o�o�oqo *<N`�o�� ����m��&� 8�J�\�n�������� ȏڏ�{��"�4�F� X�j���|�����ğ֟ ������0�B�T�f� x��������ү��� ���,�>�P�b�t��� �����ο��ϟ���������:�L�^�6πϒ�l�,~���v������ ��A�(�e�w�^ߛ� �߿��߸������+� �O�6�s�Z���� �������O'�9�K� ]�o������������� ������5GYk }������ �1CUgy� �,����	// �?/Q/c/u/�/�/(/ �/�/�/�/??)?�/ M?_?q?�?�?�?6?�? �?�?OO%O�?IO[O mOO�O�O�ODO�O�O �O_!_3_�OW_i_{_ �_�_�_@_�_�_�_o o/oAo�eowo�o�o �o�o�_�o�o+ =O�os���� �\���'�9�K� �o���������ɏۏ j����#�5�G�Y�� }�������şןf��� ��1�C�U�g����� ������ӯ�t�	�� -�?�Q�c�򯇿���� ��Ͽ�󿂿�)�;� M�_�q� ϕϧϹ��� ����~��%�7�I�[�hm��V`���V`����߼����������,��3��� W�>�{��t����� �������/�A�(�e� L���������������  =$asRo ������ � '9K]o�� ������#/5/ G/Y/k/}//�/�/�/ �/�/�/?�/1?C?U? g?y?�??�?�?�?�? �?	O�?-O?OQOcOuO �O�O(O�O�O�O�O_ _�O;_M___q_�_�_ $_�_�_�_�_oo%o �_Io[omoo�o�o2o �o�o�o�o!�oE Wi{����� ����/�6S�e� w���������N���� ��+�=�̏a�s��� ������J�ߟ��� '�9�K�ڟo������� ��ɯX�����#�5� G�֯k�}�������ſ ׿f�����1�C�U� �yϋϝϯ�����b� ��	��-�?�Q�c��� �ߙ߽߫�����p�� �)�;�M�_��߃��@����������p�����p�����,�>��`�r�L�, ^��V���������� !EW>{b� ������/ S:w�p�� ���//+/=/O/ a/p�/�/�/�/�/�/ �/�/?'?9?K?]?o? �/�?�?�?�?�?�?|? O#O5OGOYOkO}OO �O�O�O�O�O�O�O_ 1_C_U_g_y__�_�_ �_�_�_�_	o�_-o?o Qocouo�oo�o�o�o �o�o�o);M_ q��$���� ���7�I�[�m�� �� ���Ǐُ���� !��E�W�i�{����� ��ß՟�����/� ��S�e�w�������<� ѯ�����+���O� a�s���������J�߿ ���'�9�ȿ]�o� �ϓϥϷ�F������� �#�5�G���k�}ߏ� �߳���T������� 1�C���g�y���� ����b���	��-�?� Q���u����������� ^���);M_�6�a�6�����������,��7 [mT�x��� ��/!//E/,/i/ {/b/�/�/�/�/�/�/ �/??A?S?2�w?�? �?�?�?�?���?OO +O=OOOaO�?�O�O�O �O�O�OnO__'_9_ K_]_�O�_�_�_�_�_ �_�_|_o#o5oGoYo ko�_�o�o�o�o�o�o xo1CUgy ������� �-�?�Q�c�u���� ����Ϗ�����)� ;�M�_�q�������� ˟ݟ����%�7�I� [�m����h?��ǯٯ �����3�E�W�i� {�����.�ÿտ��� �Ϭ�A�S�e�wω� ��*Ͽ��������� +ߺ�O�a�s߅ߗߩ� 8���������'�� K�]�o�����F� �������#�5���Y� k�}�������B����� ��1C��gy ����P��	 -?�cu��Ы������>������/ -�@/R/,&,>?�/ 6?�/�/�/�/�/?�/ %?7??[?B??�?x? �?�?�?�?�?O�?3O OWOiOPO�OtO�O�O ���O�O__/_A_P e_w_�_�_�_�_�_`_ �_oo+o=oOo�_so �o�o�o�o�o\o�o '9K]�o�� ����j��#� 5�G�Y��}������� ŏ׏�x���1�C� U�g�����������ӟ �t�	��-�?�Q�c� u��������ϯ�� ���)�;�M�_�q� � ������˿ݿ���O %�7�I�[�m�φ��� ����������ߞ�3� E�W�i�{ߍ�߱��� ��������/�A�S� e�w���*������ ������=�O�a�s� ����&��������� '��K]o�� �4����# �GYk}��� B���//1/� U/g/y/�/�/�/>/�/��/�/	??-???��A;�����j?|?�=f?�?�?�6,�O�?�OO�?;OMO 4OqOXO�O�O�O�O�O �O_�O%__I_[_B_ _f_�_�_�_�_�_�_ �_!o3o�Woio{o�o �o�o�/�o�o�o /A�oew��� �N����+�=� �a�s���������͏ \����'�9�K�ڏ o���������ɟX�� ���#�5�G�Y��}� ������ůׯf���� �1�C�U��y����� ����ӿ�t�	��-� ?�Q�c��ϙϫϽ� ����p���)�;�M� _�q�Ho�ߧ߹����� �����%�7�I�[�m� ������������ ��!�3�E�W�i�{�
� �������������� /ASew�� �����+= Oas��&�� ��//�9/K/]/ o/�/�/"/�/�/�/�/ �/?#?�/G?Y?k?}? �?�?0?�?�?�?�?O O�?COUOgOyO�O�O��O���K�������O�O�M�O _2_V,oc_o�_ n_�_�_�_�_�_oo �_;o"o_oqoXo�o|o �o�o�o�o�o�o7 I0mT����� ����!�0OE�W� i�{�������@�Տ� ����/���S�e�w� ������<�џ���� �+�=�̟a�s����� ����J�߯���'� 9�ȯ]�o��������� ɿX�����#�5�G� ֿk�}Ϗϡϳ���T� ������1�C�U��� yߋߝ߯�����b��� 	��-�?�Q���u�� ���������� )�;�M�_�f������ ��������~�%7 I[m������ ��z!3EW i{
����� ��///A/S/e/w/ /�/�/�/�/�/�/? �/+?=?O?a?s?�?? �?�?�?�?�?O�?'O 9OKO]OoO�O�O"O�O �O�O�O�O_�O5_G_ Y_k_}_�__�_�_�_��_�_oo��!k}������Jo@\onmFo�o�o|f,� �o��o�o-Q 8u�n���� ���)�;�"�_�F� ��j�������ݏď� ���7�I�[�m���� �_��ǟٟ����!� ��E�W�i�{�����.� ïկ�������A� S�e�w�������<�ѿ �����+Ϻ�O�a� sυϗϩ�8������� ��'�9���]�o߁� �ߥ߷�F�������� #�5���Y�k�}��� ����T�������1� C���g�y��������� P�����	-?Q (�u������� �);M_� ������l/ /%/7/I/[/�/�/ �/�/�/�/�/z/?!? 3?E?W?i?�/�?�?�? �?�?�?v?OO/OAO SOeOwOO�O�O�O�O �O�O�O_+_=_O_a_ s__�_�_�_�_�_�_ o�_'o9oKo]ooo�o o�o�o�o�o�o�o�o�#5GYk}���$UI_INUS�ER  �����q� � ��_ME�NHIST 1D��u  �( �p��.�/SOFTPAR�T/GENLIN�K?curren�t=editpa�ge,LABWE?LD_2,1�H��Z�l�z)	��MA�IN5�ŏ׏��� �'���menu'�71��G�Y�k�}��q(�#�95,18��Ο��������?,148,2�R��d�v����)�,15�46�ԯ���
�p/���AB_/�5�^� p����#�5�G�4��������p�(��3�E�W�i�{ύϟ�  /����������߭� B�T�f�xߊߜ�+��� ��������,��P� b�t����9����� ����(���L�^�p� ��������G�����  $6!�Zl~� �������  2D�hz��� �Q��
//./@/ R/�v/�/�/�/�/�/ _/�/??*?<?N?�/ r?�?�?�?�?�?�?m? OO&O8OJO\OGeO �O�O�O�O�O�O�?_ "_4_F_X_j_�O�_�_ �_�_�_�_w_�_o0o BoTofoxoo�o�o�o �o�o�o�o,>P bt����� ���(�:�L�^�p� ��mO���ʏ܏� � ��6�H�Z�l�~��� ���Ɵ؟���� � ��D�V�h�z�����-� ¯ԯ���
����@� R�d�v�������;�п �����*Ϲ�N�`��rτϖϨϓ��$U�I_PANEDA�TA 1F������  �	�}  fr�h/gui��de�v0.stm ?�_width=0�&_height�=10	���ice�=TP&_lin�es=15&_c�olumns=4�	�font=24�&_page=w�hole���ϑ�)�  rimX߁�  ���ߪ߼������� Y��(��L�3�p�� i��������� ����$�6��Z���� ��  z� N�>�ߗ������� ����D���9K] o�������� �#
G.k} d������n�&��6;/M/_/q/ �/�/��/,�/�/? ?%?7?�/[?m?T?�? x?�?�?�?�?�?O�? 3OEO,OiOPO�O�O/ $/�O�O�O__/_�O S_�/w_�_�_�_�_�_ �_J_o�_+ooOoao Ho�olo�o�o�o�o�o �o9�O�Oo� ������r_ #�5�G�Y�k�}���� ��ŏ׏������1� �U�<�y���r����� ӟFX��-�?�Q� c�u�ȟ�����ϯ� ���~�;�M�4�q� X�������˿���ֿ �%��I�0�m��� ������������b� 3ߦ�W�i�{ߍߟ߱� ��*��������/�A� (�e�L������ ��������Ϟ�O�a� s�������������R� '9K]��� h������ �5YkR�v�&�8�}���/!/3/E/W/)�|/�� k/�/�/�/�/�/?i/ &??J?1?C?�?g?�? �?�?�?�?�?�?"O4O�OXO��B�<��$U�I_POSTYP�E  B�?� 	 dO�O��BQUICKME/N  �K�O�O��@RESTORE� 1GB�?  �KO��!5_BS0_��m`_�_ �_�_�_�_t_�_oo +o=o�_aoso�o�o�o T_�o�o�oLo'9 K] ����� �~��#�5�G��o T�f�x����ŏ׏� �����1�C�U�g�
� ��������ӟ~���� �v�(�Q�c�u����� <���ϯ�����)� ;�M�_�q��~����� �ݿ���%�ȿI� [�m�ϑϣ�F������������GSCRE��@?�Muw1sc*Pu2J�U3J�4J�5J�6J��7J�8J�'�TAT��M� �CB��JUGSER,�1�C�T+ЦL�ksT���4��5*��6��7��8�ъ@�NDO_CFG �H�K���@PD������N�one�B��_IN_FO 1IB�q��@0%ߌ���z� ����������'�
� K�.�o���d�����������L^�OFFSEOT L�Iu��� ��#P��,>Pb� ������ (UL^���@���O��/
/�:/��UFRAME�  ��.�[�R�TOL_ABRT8^/Y�v"ENB/p(?GRP 1MY�ACz  A��# �!3��/�/�/	??-???Q;r&�@U�(3�+?MSK  �%q�ڎ+N[!%i��%x��?�%_EVN~ b�4-��6�2N
�
 h3�UE�V~ !td:\�event_usger\�?B@C7GOd/��F|L:ASP@A�EGspotwe{ldwM!C6�O}O�O*P�4!�?VO_ I_�G�1_8_&_|_�_ \_n_�_�_o�_�_�_ So�_wo"o4ojo�o�o �o�o�o�o+O�o �0��fx������zFWRKg 2O��&!8�y��� g������ ��ӏ�.�	�R�d�?� ����u���П�������*�<��M�r�����$VARS_CO�NFI"�P
 F�P�����CMRv�"2V
�9��	4ೠ��1:� SC130EFG2 *���ę�Y��x�0�5��3�?�a0@a0pU0�N�� )/h�r� �ȓ���ҿ��Ϳ��k�-O5A���7���� B��� R���V�޿wϾ���j� �Ϫ���������=� ���s�^�pߩ�\���|�ߓ�IA_WOQ��Wi��v,		��F�(�6�G�P ��I��H��RTWINURL ?&I���ߎ������������SION�TMOUO �� �BXS۳��S۵@�! �FR:\�\DA�TA�O  ��� MCA�LOG�N�   UD1�A�EXr���' B@ �����`����������x �� n6  ������6��  =���M��J ��g�TRACIN��\�Bd��pMQ����ңY&K (�ѝ	��� ��%[I m���������_GE)�Z&K�`
��
� 
�?"'��RE,�[�)�����LEX $\���1�-e��VMPHA�SE  &E��N���RTD_FILTER 2]&K �1��_� ?? $?6?H?Z?l?~?�?�? ��/�?�?�?OO*O�<ONO`OrO��SHI�FTMENU 1�^�
 <��%���O����O�O_ �O�OC__,_y_P_b_ �_�_�_�_�_�_�_-o�o	LIVE/�SNA��%vs�fliv�.?o�}� SETU��bbmenuxo}oo �o�o#�E)�_k�HkMO)�`.�z��KZDta\/
�<���P�$WAIT?DINEND��|!rvvOK  �ȑ|��S��yTI]M����|G} ��0�������xRELE�!@�v�vs��xq_ACT�U`?��x_J� b��%�o@����ORDIS����vp�V_AXSR|�2�cYyw�D(|�Ӡ_I�R  �&t�  7
ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v���ϚϬϾ�NXVR�y!d7~�$ZA�BC�1eY{ 	,� ��2����Oq��VSPT f7}\�r{�
�j�o����j�ߣ�B�DCS�CH{ g�d���I-PRrhY�6��H�Z�l���MPCF__G 1i��05X׫�q�MP�j�66 p5������<�0  ��ܳL?y?�O���  �����3\�K4��+�+�&�'���Dd�8C�����?�?�=ۄ�4 �{���&�8�J�1V���z�?����������/��� �d��ð�XD̿73����W���3�FX?��� ����~�����P�A0��C�Ą�{ k��W_CYLIND��!l�� й�? ,(  *����Ӧ��/�   =/O/a.��/��/ �/�/�/!/??&?i/ J?�/�/�?g?�?�?�/0�?�?O��2md� ġ�7OGLj��pO[O�O��'O�O�ז��AA�wSPHE_RE 2n��>? _�?_P_7_t_�?�O �_�_8?�__e_o�_ :o!o�_po�o�_�_�o +o�o�o�oYo6HlZ��ZZކ �ʆ