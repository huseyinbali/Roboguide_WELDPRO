��   �A��*SYST�EM*��V9.1�0214 8/�21/2020 A   �����
�WVAMP�_T   �$X1  �$X2AY@���/FC5  �$2ENBA $DT  / �_R2 d E�NABLEDnSCHD_NUMA �SCFG5�� $GROU�P�$z ACCE�L@�G$MA?X_FREQ�2 �L�DWEL�D�EBUG�PRE;WSOUT��PULSEAS�HIFt 7TYP�4$USE_A�EF} 4$GD=O�  f0� r?�NpW�EAVE_TSK� �V�_GP��SUPPORT�_CFnCNVT_DONE p �}k}GRP #2r�� _� ��$� TIME1�o$2'EXT�� (1#&(MODE�_SW�CO3 S�WIT � TPH�AX6  4 �� ECC$�T�ERMNnPE�AKno!AL � \ � �!I֑$�!N_VSTAR�#!r"ؾ�"�%�CY�CL42 
�S� Tv"b $�CUR_REL_�� �!3WPR5� � 
$CEN� _RI3RADkIU�XI�z ] ZIMUT�i!$ELEVAOTIONg5� N��CONTINUO�e2q �MEXAC=PE� x�6 � H~ �UEN�CYA�ITUD<4�2RIGHC�2�LEBL_ANG�1 �OTF_�� 	�  1$3A�bET���n3C!$O;RGjHFBKjH���P��C��DLD%W�HR�E�_�3�B �C��D�B�C�@�D�A�CCHG�G	Q�F	Q8�F	Q�FINC�G=Q �F=Q�F=Q�F�AVCPYC� _T�\#�Y�~P#�@SY��H)@�UPD"0n��$$CLASS  ����Q���8 �P�PVERS��1�W  ���QIRTU�AL�_�Q0 2~�X�  ��{?��@�  Ha Dae�TWoio{o�o�o�`)dN 2 3k� Hf��uHe@O�Hi�oNc)a� � e� E`��i ��Ca��d �`z����=�����4s ����jpYq8��w�r��
|�{ at��ujp`��i.�5t8q�q2�b�t���
�<q`����� Ca����̏ҏ�����)a�  23k
{TDaSI�L8� �������h�?m�'����l�D� ����Ca��l����k�� � �2�D�V�h�z��l�FIGURE 8��o�v�Ha l�f��������M� (�H��󈯎�����Ŀ�ֿ�TCIR1��Pd�}�0�~�`h�z�D�Z�l���0� v˜�~����� ��$�n�jN� 2��4q�Ȓ���@��ʖD� M`g����������	��-�?�Q�c�u�`�� �q� �5)�ᐟN`���� ������˟���M�_��q������������k�Triangle��z�h߾�M ��Ɵ�ύ����`��/ L� &��g�n� ��	//-/?/Q/c/ u/�}DVhz��/ �/��9?K?]?o?�? �?�?�?�?��Lu�� Oe��O2ODOVOhO zO�O�O�O�O�O�O�O 
__.[�?._O"O�_ �_�_�_�_�_�_oo�&o8oJo\ono�mSC�HEXTENB � =��ctSTA�TE 2�k �|o�o�o �gWPR 7�6�L}�D�-�_OTF 		8��@)0�q�q�0��v)��uAȫs�u�@�  <#�
��?����mu_GP; 2w| ��� d�v����я㏡+