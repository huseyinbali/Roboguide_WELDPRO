��   ��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	��/GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1  	��CLo�: � �A�X{  $PS_��TI���TI�ME �J� _gCMD��"FB��VA �&CL_OV��� FRMZ�$DmEDX�$NA� �%�CURL��W���TC�K�%�FMSV��M_LIF 	��'83:c$�-9_09:_��=�%3�d6W� �"�PCC�OM��FB� M��0�MAL_�E�CI�P:!o"DTYkR_|"�5:#N�1END�4��^o1 l5M��P PL� W ��  $STA:#T�RQ_M��� K$NiFS� uHYsJ� *hGI�JI�JI�E#�3AZCaB�A����$�ASS> �S���A�����@�VERSI� �G�  �~QIRTUAL�O�QS 1X� ��� 	 ��x_c_�_�_�_ �_�_�_�_ojP5f Be&m Q^oLo��2P�A� �YUV��XHso�ooql�o�o�o$�kW]rF ������d��x����=L���f8�?�9���@�Y� ~�������Ə؏���`� �2�D�� 1U�o�}�g����D  2 �Ο�����(�:�L�^�p���<������ ��Я�����*�<�8N�`��j	 (��� �����ܿǿ ���� 6�!�Z�E�~�iϢύ������$4 1�N\���L�:��L�l�K�f��O(LP�K�K�Ո��A�+@�xr@w��h<8	�<�k_(<$�4��@L� \ߵ��ϕ߀߹�T�f� ���ߤ�1��U�@��y���Wzr�W��t���� ���p���l�����1�C���%��345?678901c�k� ��񍟨��������� ��`�"4��
�� d���v��� �J�*N<r �����\� //8/��q/�� �/"/�/�/�/�/T/%? 7?�/�/j?X?�?|?�? �??�?>?P?�?�?O TOBOxO�?�?�OOO �ObO_�O_>_�Oe_ w_�O,_�_�_�_�_�_ oZ_+o~_�_
o�_^o �o�o�oo o�oDoVo $�oH6X~�o� �
l����2� D��k���J���� ԏ��N�`�1����� d�⏈�v������� ��J���*��N�<�r� ��ڟ�������\�ޯ ��8�����q�į֯ ��"�ȿ��ؿ��T�%� 7ϊ��j�Xώ�|ϲ� �����>�P��Ϝ�� T�B�xߊۙ��ϱ�ݎ,�!X����U���$PLCL_GR�P 1o��� p(�?�  "�4�,�W�(�{� f������������ ��A�(�2�t�