��   ?Q�A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N  &S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  ���!IRTU�AL�/�!;LDU�IMT  ���� ���4MAX�DRI� ��5
�4.1 �%� � d%	 ��}? i?�?���" ���?�?�? O�? �?6O�?3OlOO-O�O QO�OuO�O�O_�O2_ �O�Oh__�_;_M_�_ �_�_�_�_�_.o�_Ro ooMo�oIo�omoo �o�o*�o` �3E�i��� �&��J������� }���e�w�쏛���� я�X�C�|�+�=��� a�֟����џ�͟B� ��x�'�����]��� 䯓����ɯ>��;� t�#�5���Y�ο}��� ���:����p�� ��C�UϏ����� ߯� ��6���Z�	��Uߢ� Q���u߇��߫� �2� ���h���;�M��� q������.���R� ����������m�� ��������`K �3E�i��� �&�J��/ ��e���/� �F/�C/|/+/=/�/ a/�/�/�/??	?B? �/?x?'?�?K?]?�? �?�?O�?�?>O�?bO O#O]O�OYO�O}O�O _�O(_:_�O#_p__ �_C_U_�_y_�_ o�_ �_6o�_Zo	oo�o�o �o�ouo�o�o�o �o �ohS�;M� q����.��R� ����7�����m��� 􏣏�ǏُN���K� ��3�E���i�ޟ���� �&��J������/� ��S�e����ׯ��� ѯF���j��+�e��� a�ֿ����ϻ�0�B� �+�x�'Ϝ�K�]��� ����߷���>���b� �#ߘߪߕ���}ߏ� ��(�����#�p�[� ��C�U���y����� ��6���Z�	����?� ����u������� �� ��VS�;M� q���.R �7�[m� ��/��N/�r/ !/3/m/�/i/�/�/�/ ?�/8?J?�/3?�?/? �?S?e?�?�?�?O�? �?FO�?jOO+O�O�O �O�O�O�O_�O0_�O �O+_x_c_�_K_]_�_ �_�_�_�_�_>o�_bo o#o�oGo�o�o}o�o �o(�o�o^[ �CU�y��� $�6�!�Z�	����?� ��c�u������ �Ϗ �V��z�)�;�u� q�柕����˟@�R� �;���7���[�m�� ��߯�ǯٯN���r� !�3�������޿���� �ÿ8����3π�k� ��S�e��ω��ϭϿ����F���j��+�
S�end Even�ts�S�SEND�EVNT��Q��އ� %	��Da�ta�߶�DATA�������%��S�ysVar;��S�YSVw����O�%�Get�x�G�ET+����%�Request �Menu���RE�QMENU?���� �]ߞ�Y���}�+��� ��.��d� 7I�m���� *�N���� �i{��/�� /\/G/�///A/�/e/ �/�/�/�/"?�/F?�/ ?|?+?�?�?a?�?�? �?O�?�?BO�??OxO 'O9O�O]O�O�O�O_ __>_�O�Ot_#_�_ G_Y_�_�_�_o�_�_ :o�_^oooYo�oUo �oyo�o �o$6�o l�?Q�u ����2��V�� �������q����� ���ˏݏ�d�O��� 7�I���m�⟑���ݟ *�ٟN������3��� ��i���𯟯�ïկ J���G���/�A���e� ڿ�����"��F��� �|�+Ϡ�O�aϛ��� ��߻���B���f�߀'�a߮�]��߁ߓ���$MACRO_M�AXX�������Ж�SO�PENBL ���2��ݐ���_���"�PDIM3SK�2�<�w��SU���TPDS?BEX  K��U)�2�����-�