��   K�A��*SYST�EM*��V9.1�0214 8/�21/2020 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_���$$�CLASS  O�����D���DVERSIO�N  ��/IRTU�AL-9LOO�R G��DD<x$?�������k,  1 <DwX< y�����C�����	/��Z�Zm//�/�_/�/�/�/$ ��/�/	?';�$MNeU>A\"�  �<�������'�?h0�c11�m�'��&�'��5!C���l����Ý����0��NV��~��¹�?�˼N������J���·�?~��C�"�CZNÚ��:5/�?�� �?�?#O	O+OYO?OqO �OuO�O�O�O�O�O_��O%_C_)_97NUM  ����w92�TOOLC?\ �
Y7?O�_Ry3\�N�TPﳗ�P�R��.���P©� &�?�5C��o7_Y_ 	o1_o?o%o7oYo�o mo�o�o�o�o�o�o�o ;!CqWy� ����sV�Q�Vy �[