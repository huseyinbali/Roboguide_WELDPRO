��  	G��A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� ���PCOUPLE�,   $�!PPV1CES C G1�!IME A> �1�	 � $S�OFT�T_ID�BTOTAL_EeQ� Q1]@NO`B�U SPI_IND�E]uEXBSCR�EEN_�4BSIG�0O%KW@�PK_FI0�	$THKY�GP�ANEhD � D_UMMY1d�D��!U4 Q!RG1R��
 � $TIT1d ��� 7T@d7T� 7TP7T55VU65V75V85V95W05W>W�A7URWQ7U�fW1pW1zW1�W1��W 6P!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2� � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1�0UT�OB U��0 9DEVI%C4ST3@�� P@�13��`BQdf"VA�L�#ISP_UN9I�#p_DOv7IyFR_F�@K%D1�3�;A�c�C_W�A?t�a�zOFF_�@N�DEL�xL�F0q�A�qr?q�p�C?�`�A�E1�C#�s�ATB�t�?
�WELDH2/0 =s�qn"QING�0$��QA7PD2�4%$AS$d3�BEl�P�_��B�UCC_AS�BFwAIL��DSB��gFAL0��ABN@��NRDY���`���z��YN��SCH���pDE���yp���������|�STK`>���	���	�NOj� ?�ڂL��d�U* G� ��9 ���������߇�ƗƗ��ԘS_FbәE��F�ƗSSŘ2��P�1 �ON�F��HOU�D�MI:�1D�SEC`B�2yi �HEK0~���GAP������I�� � GTH���0D_ȡ����T= ��� ��
��p}�9!K���9!ƗUN14��5���#MO� �sE 	� [M�s��t�REV�B����!�XI� g�R � � OD}`��i�`M�m�����/�"��� ŵ��eaX�@Dd �p E RD_E����$FSSB��&W`KB!�E2uAG� J��  "��S��� V�t:5`�QC=;m��a_EDu � � C2�f��S�pa�l �t$O�P�@QB�q��_OyK"�آTP_C� ���da�U �`LAC�m�^��J�� FqCOMM� K�D��р@�p���OR�BIG�ALLOW� �(K\��@VAR�w�d!�A}!�BL8[@S � ,KJq��H`S�pZ@M_Ox]�՗�CFd7 X�0GR@�z�M�NFLI���;@Uɠ�84�"� �SWI�&"AX_ANo`����9��G�� �0WARN!Mxp�d4�%`L�Tb\;�� COR-r�FLTRY�TRA�T T�`� $ACC@�TB� ��r$ORI�.&�;RT�`_SFg WCHGV0I���QT��PA�I��T��e`5��� �� �#@a"��HD)RՃ7�2�BJ; �CTO�I�3J�4J�5J�U6J�7J�8J�9��xȰx@�2 @� TRQ��$%f�������_U��������COc <� ����
�3�2��LLEC��o�MULTIV4�"fѱAv
2FS�ILD��
1;�Oz@T_1b � 4� STY 2�bv�=��)2_�p�:��� |9 $�.pڰx�I`�L* �TOF �sE�	EXT3ء�B3��22�0��@�	1b.'.�}!9�
���  �"�� /%�a�g�?s���!��;AآM��`Q  �T}RE� " L�0��	�`��pA�$JOB��E����$;IG� # d�,/ >/P(���#��ނ_MORc$ et�F͠�CNG�AŠTBA �6c� :/�9��0�19@�G;P/pH5���`A�%L����Bq�1��&rJ��_R�������;J@��8�<J� D 81��9Q��2�@���;�Rd&� P
	�rG�R�`�HANC?$LG w��a2q�͠�Z�/�P�
0�2�R��Li�a�D��)�CDB`f�CRA�c�CAZ�`��HELT��F+CT<�.�F"�`R�M#@�AI([O(X ����
1�Rw�w �3/�S���1��5�M�P�����HK&A�ES_SH�Q�W
��N0S��Z����_'  v@I#��Aq�Rc(��STD�_C�t�Q�3"U�ST�U��)kT�IT�a~Ф	%�1I-Oy���@_Up�q���* \����UpO�Rzs`b��}�~p�`O,~@N�SYR�G`�q �eUp�Љ�� ���L�BPXWOR�K��+��$SKد�<�p1DB�TR��p , ��0A`���c�B��W�DJDS _Cdд�sDPwPLzq�ё�s��DM�<wY����2��2H�9N�p� Eb�A2��-�bHaPRi�M��

�D�� ��.� q��1$�[$Z���L�y/�&������0���w�P� 1���tENE��� 12��s~pREv��r3H $C��o.$L`�/$�s8���tw�INEV�a3_D}�m�RO3��� I;�~!�`�:���?RETURN��2�MMRj"U琋�C�ʠNEWMA`#�S�IGN��AJ@#�L�A<�!�&P0$=Po 1$P�@�24�M�;�O�� S���a�o��v�Q�V�GO_AWT #�`��@`ъQW�DC,)�o�CY� 4'"��1�(����Ĕ2��2�̖Na���C�4��D�EVI�� 5 oP $��RBUÖ�PI̗P��3�IG_BY�;�J�T�1��HNDG�q6# Hv�c&�E�g� ���#�㗣͖�`���L�7w��`�Ѭ�3FBڬ(�FE������͔��@�ܱ8� p�МQ��@�MCS4��Ƞ�dH����RHPW�F��5:�J n���S�LAV.�9�INP��J��Ш����_:P +B�S6@�`�� B�� 1�FI(b��	��5Oa�Q'OaW	�NTV��V��SKI�CTE*�@��b�]�&�QJ_S�R_����SAFv�5���_S}V2EXCLU*v`-�D~`L����Y�{�HI_V<RP�RPPLY4px�p��u�۶��_ML��v`$VRFY_ts��M�IOC\��%C_>PS�T�]�O�/���LSр��nt4�Fqy�͓� �`P��en⯐K�AUNF����͕���ZqCHD�$������ �AF� CPU#��T�Fqĳ?Pס ;�4��`T��c�� ���N�� <$��8@TЀ�� ��g�óSGN=�0
$U0������Б� �*0e �b��b��ANNUN�����͕U0�4v`'�w ����>PX�����EF�`I�>��$F��&dO0OT��nt��prTqh��kq)�M��NI�r!?'"|�G~�Aޱ���DAYecLOAD��ctu�os5v�EF_F_AXIɢ@4��Yq�SO���s�`_�RTRQ�A D�y�Q� Qt` BE���� @�P��WP  ��AMuPC@E�� B��XT]2Xl�8FDUt�8E��bCAB��C8�*�NSj0ID�!WRBU�A:P�V%�V_T  �@��DI%0cD� �1$V�SE�T �2]3�1�o�
��]2f�1E_��lVEP	0SWAQ�0�� 3  AN0��O�HqPPAmI	RAa]2B�`�n�� ���S��@�@�%�� C�P ���RQDW�MS��P%AXt/lLIFEp�. uq:"�NA!M2J%��?#M2C�����C�P��N0�$ǁ�&��OV��V&sHE��]2SUP�!��:"p_�$��y!�_:3�%���'Z�*W��*�Q�'S�ሢ�RX�Z�@�qY2=8C"��T�`��	N?�*��J%Q �_�@� J�I@�TE =`�CACHt���3SIZp&� ��%��NZ�UFFI� ��p��ct��os6�wry�M�P%DF 8���KEYIMAG�TM���C#A��F���Ɓx�OCVIE$K�aG�R�@LCĐ�^ �?� 	#�D?Pj�4H b�STo�!�B�ГDTp�D����D��@EMAIL��𽀣����FAU�L�rI�R���cPC#OU�PFAJ�TO��Q?J< $�C5��ST � IT��BU�F�7 ��7
�4`*`� B*T5�C�����BAcPSAVuU7R @\2:�U�W����P|T5�R�L��_*P[U��F�YOT���`��P2�0\p�Z?��WAXec+�b=�X*P�éS_GA#�
� YN_���K� <� D0�!p����M�� T��Ffƀ$݀��DI �!E�`O�P��aL����	GKQF�&�㌁�a��8����	�M�\��aL�C�SC_��K���`���d��RA�e�H��aDSP3F�bPC*{IM�S!sGq��a�� U�g� ��"��@I�PD��c{0 tTH�[0��r��T��!sH9S�csBSCQ�j0*�Vְ�z�p!c�tf���NV��G ��t[0$v*PFAB`ds}`�aǁSC�&��cM�ER��bqFBCM�P���`ET�� mNBFU� DUP0���22��CDy�pl�P�CG�ЀNO��
��O �����R��PN�Cj�υ�R�@b�A���P��P/H *ρL۰�� ��QL����o�B��� @�j�@���@���@��1*@�7=�8=�9=�A T?�I�1V�1c�1p�U1}�1��1��1���1��2��2I�V�2�c�2p�2}�2��2���2��2��3��3RI�3V�c�3p�3}�U3��3��3��3��94���AEXT���QTb��Y`m&Y`:�d`t���"�FDR�/RT
PV���Rp:"ɱ�r:"REM#9FU�OVM�cﵽA��TROV��D�T�P�MX'�INp��� ��IND6�B
bȎ`B`W`G*a �!��@J%0D!��RIV�n"GE[AR�aIO'K�lN}`����%(L�?@|� mZ_MCM50n:!��F� UR{��S ,́MQ?� � \p?4�@?4�Et�<�H�gQ�X���T�0�Pa�� RI����8RE�TUP2_ U ��6STD�px5T�T��LѢלչ�7RB;ACNbV T��7R
�d)�j%<��x`�IFI�x`X�)�A ���PTM�AFLU=I~DW �� `H PUR�`Q�"�R�aP�p-P�$ Iܴ$p�]S$�?x|�J�`sCO�P�SVRTl�>G�x$SHO#���CASS�p�Qp%�p��BG_���V����c���p���}�FOR�C�B -�DATAZ��X�BFU�1�b�"�2�a��/�[0��Y� |r�NAV`S�p����S�B~n#$VISI��6vbSCdSEZм�V��O���B��I� ��$PO�t�I��FM�R2��Z  Ȳ���ɱ�`��ͷ��@������@�_��9��$IT_ᛄ�"M�Ʋ���DGC{LF�DGDY�LDLѐ�5R&��J$��0��~E[G@;	� T�FS�PD\� Pz��cB`$GEX_.1`���"3P5P�9G�q��] �L�x��SW^UO�DEBcUG���GR�к4@U?�BKUJ�O�1� O PO@ ��j���M��gLOOc�SMK �E�R�AT�� _E �^ 7@�� �/TERM %_)&�0'ORI�a% `)%��GSM_�`��% a)%h��h(bB)UPUB�c� -S��Q^p�7#� _��G�*^� ELTO�q�b�FIG�2�aЛ�,@N$�$`$UFR�b$À�!0��fV OT7�TA�p�ɰ13NST�`PA�T�q�0G2PTHJ�n���E�@�R���"ART�P�%�@�Q�B�a�REL�:9aSHF�T�r�aM1{8_��R(w���f& q $�'�0�bvʰ��\s9bSH�I�0sU9� �QAYLOvp2aHa1�]���M1B�ׅ�pERV H�Af��8l�-7�`�2`��sE��RC\�ׅASYM{aׅ�a#WJ�'l�h�El�w1�If◁U�D�`Ha{5� gF�5PZs5@
��6kOR�`M��Tw!��d��L00�1a�HO���e a�S1��OC�!���$OP0���a.���䱩���`䰚PR�9aOYU�sM3eV�RK5��U�X�1��e$PW�R��IM�UIBR_��Sp4r�g `3�aUD�lӳ3SV	�eQ�df���$H�e!f`AWDDR��H!GO2�atamaj��`���g Hz�SE���壬e`�ec��ep�SE?̐�i�HS����h3 $��P_Dq������bPRM_R��|!HTTP_H��i (��OBJ؊�mb��$��LE�>3cP)q�j � �|�b�AB_c�T�#{rSYP�s@�KR�LiHITCOU �t���P��P{r��l�0��P�PSSg�;��JQUERY_F�LA�!b�B_WE�BSOC���HW����!�k�`�@IONCPUdr�O:� �qH�Q��dR��dR�p���IOLN��l� 8z�R��d�$�SL��$INP7UT_!$�P���P��  }�SL]A� m�����مՄ�C���B�aIO^pF_AS�n�Ї$L��Ow���1 ��"b�!I������@�HY��X�1�n��U;OP�o `�v����F�H�F�O����PP &c�P����O�ǒ��h�ru�M�A6�p l6� CTA0BVpA��T�I���E&P ��0PmS�BU IDC  �r��?��P>�|!�:�&?0qЂ��+��⩀N�� ���IR�CAڰ�� r ��myԀCY�`EA@�͡��ҬF�&c��k�Rg0�AA��ADA�Y_G�B�NTVA�E�V�.�Ȃk5:�.�S3CA*@.�CL��G�"���G���6�sr���Xl2����N_�PC���G��7�tЂ�S ޱ��JrG�>�p"�� 2se����6��u���Jr�LABp?13� 9�UNI�9'�Q ITY���$xe�R���vЂM��R_URLT��$AL��EN�n�s�tg �TrqT_Uk�� �J9�6�w X �����E��9�R����"] A�Ӂ��Jv���#FL9k���
Ӻ�
�UJR��x �mpFA�7��7<ҽD{�$J7��O^�B$J8g�7PH!�p҂�78�c�8���f�APHI� Q�qӶ�D+J7J8�����L_KEd� � �Kt�LM��� y <��X�R�G�ţWATCH_VA��5@~�Fv_FIELDhey��L�ҁ�z R 51V>@¦K�CT��W�
�r�:�LG��{�� !��LG_SIZut���� �����FD��I������ ��" ���S����  ������" ��A8�� ��_CM#3`���g�-F�An�����r�T(���2�ိ�� ��������I��������" ����RyS�\0  (�SLN[р|���p �@ڂ��,��s:rYPLC9DAU_�EApt�|Tuk GqH}R�a �BOO�a?}� C7� `�IT�s�03�RE��SCR��s8��DI2�S0RGI"$D���+��TH�t �S[s�W�� �N+�JGMTMgNCH� �FN��bWK}��{UF���0�FWD�HL.�STP�V�Q X�� �RS�HP�(�C�4��B+�=P0T)Uq�/��>�a�@��Gm�0PO��'���i�sOC�EX'�TUI{I��ĳɠ��4	1�E3yd��0G���	�c���0�NO6AcNA ��QD�AI9�8ttt��EDCS��c��3�c�2O�8O�7S���2�8S�8IGN��G���zm��43DEOa5$LL�A��HAT��~F�u�T��$��l�B�ä���-A\aF��P��PM�p�� 1�E2�E�3�Av��!�0 �m{Qk3������?�=Q�u� ����FST��Rv Ys�R0P� $E$VC $[[�p3VFV `��$ L4�F��P[�`=�[����Q$eENp�$d%6�_ ���q�q`�� �S ��MC-� ��9�CLDP����TRQLI]���	i�TFLGR�P�a+cr�1D:�+g%�LD+ed+eORG��/!>bU�?RESERVU��d��c�d�b��S�c� � 	e/%d+e#SV 	`�	na�d}�fRCLMC�d@�o�oyw��a`�M�p���Ѕ��$DE?BUGMASI��H	�Q�uTu05�E���TQ�MFRQ~��� � ��HRS_RUہ�Q�A�T%FRE�Q��Q$%0��OVER-���o��FA��P�EFIN�%��Q�]q[��s�d�� \���q��$U��@޲?�`G�P)S�@��	�sC~ �c��W�sU��bq?�( 	v�MISC�.Ո d6�ARQ���	��TBN� 1��&1ˈAX�R��|·�EXCES�¤�Q��M���щm�����T�R��SC�@ O� H۱_�����S�����`JP�T�ċ &�i�F�I��MI�� �� �Po�^�H RCT�Ns��ȖOҚAҚ��ԐCx��u�ԐUSEDw eO�@TЏ�PX�� ��������^P)�/�+e�R� �pSZ��B_�FR�`T��\�Z_��^�CO>� PHq�K�čA�h�cuB]_��LICTB� �QUIRE=#MO���O��)�1�L�PM�Ŏ �P���r�4���b��NDK��B�Џ4+��9�Dx��GINA�DRS!M\�S��0ё�S#x��P'�PSTL��7� 4��LO̐�D�RI��EEX��A�NGk2k��ODA�u���5�=���MFm����v�I�RAp�U&�( avSUP�Uz��F �RIGG� � ��`�S'� ��SG&�T��Rn� P~�P��r��#mqPG�W�TI/��@��(�M�\�Qr� t�MD
��I)�ƕ0�q��Hϰk��DIA<���ANSW"ԨmA�!�D})HqOqR�b�`�Д ��U��VB��`k�j�9_Lp�ѕ ��@�C���Np+�����Pе� ����P��KE8I"��-$B�p��NzPND2r�a��2_TX�TXTR�A�31�%r���LO�w ���$�G�T��F�.�|�g�_�ڲR�R2���� .�W�[A�a d$OCALIĀ(�G�1:��2�@RIN���w<$R��SW0t���%sABC��D_�Jഡk���_J3:�
�1SP��r�k�P�-�3,���vP
k�\�J%sl��b�a�O.AIM%p��CS�KPj��> qs��J~��Q�����������İ_AZ�bh���E�LAg�qOCMP0ҳ��J���RT�q)�Y�1�i�G�Ȁ1��K40Y
ZWSMG� ��3tJG�PSCyL���SPH_�0�����`k���R'TER���S0��)_�0�Q�AS̊��DI�23�U��DF^P�L�WVEL	aIN8�R0&_BL�0k�.��l�J3LD�MECHPB%rP�IN� �q���|҂�2�k���sP_�� ������Ч?������DH�3഑�v@$V��R���41$v �q�r���$�a��Roӵ���H �$BEL� �w�_ACCE@4(�S'%qa ʐ_� J�q��TJ��C*�EX�RL6��&c� w'��w'.�W)�'m#�'-36�RO
�_�A!"�� 1�uu�W!_MGƺsDD!1��rFW��`��]#=5m#X"28D}E[;PPABN�'RO� EE2�A�?�	`��AOqO�X!^P��_��bSP�pC�TR�4Y}03 �a yQYN��A���6�����1Mwq�ѭr0O8 ��CINCa�̱�Z2A4˂:G��́ENC� L��k��!X"Ʉ+�IN�BI6��E���NTENT2c3_�r�CLO�r�@�pI�U��F@j��\��@ia�C��FMOSI&1y����1�s��PERCH#  k�q� .Wұ 9S���B3t��$�5$)���A�"�UL�4��t����EF��J�V�FT3RK��AY[�(� O��Q�"ecͰ/S�HB�pMOMc�˂O� �`��T�Y3��c�#̰2��DU��7�S_�BCKLSH_C �"�ewpV�p�3j��c�aB�jA��CLAL�M�D}q>`��eCH�K�����GLRT�Y���ӁD��?���_��T_UMps=vC�ps/1�Us�pLMT)�_L nt+�ywEs}�p�{rp�%�u�(�>�aA�P�trXPC�?QrXHI�۠%5=uC�MC7�/037CN_b��N6�4�t�SFE!cYV�2��wG�	��"�x��CATD~SH þ�34iF?�xaxFX�07�X�L "0PADt8B_PCu'c_�� f�"P��c&�uJA�T��a��?�'��TORQU�0/� Sii0��0R�i0��_WVe�T�U"!��#��#��I*��I��I#F尜��s�����+0VCW 0�1Wd�1%�#09���+�JRK%�j�]�u�KDB� M��u�MP��_DL!�RGRV�����#��#��H_p^㈣� תCOS�1 �LNl��(��  	�v 	�ۑE�3���b��Z�V��MY�����������THE{T0�ENK23#�β#�CBӶCB#C��AS����۔0�#�ӶSB#$�N޵GTS��1C0�� �O�_Z�B�$DUp�W£�5���DQnQ_�sjANE
���!K$t;	��±AƵ����֥�ᡇLPH��§E��S (�@�3�@�B���Q�j�(T�q���V�V� �)�V8�VE�VS�V�a�Vo�V}�V��H��*�0�(ݭ�G�E�H�S�Ha�Ho�H}�H*��O�O�O��'�UO8�OE�OS�Oa�UOo�O}�Oq�F����O�3�T��SPBALANCE_����LE;�H_ƵS�P�$���3���B�PFULC��������B��1�=UTOy_puT1T2	S"2N�a^"�@3�@7a����"N#RaT�P�O� `!��INSE9G^"�AREVX�@ΐADIF�U�1�l��1��@OB��a��dg2u��@q��?LCHWAR}2�2AB��feo�@��(
AqXsX
aP�t)8��� � 
*���L!yEROB"PCR��"l� �C�J!_�T � �x $WEIGH@i@$ӥ)��IA�@IF�1;0LAG�2�rS�2� �27BIL�OD@`�@&�STd �P��`B��1 �������
]@J"�1�  2y��D�DEBU��L� "~�MMY�9�%� N��m$i@3$D�!IQ$W $���� _C�D�O_� A�� <@�'& ���1��B���N�C�(_�@�0�"O�` ��� %\pT�@�A[qTx�O$� TICK�� T1� %3�`(0!N"P �#"PR�`�1��:5�F5� PRO�MPCE� $IRk��1p�2�P�2MAI��2A	B�5_��3� a@�R��COD,#FU�0�ID_AP�5� �{2��G_SUFF�ې ��1�152DO=7x >5�=6GR��D[3&D��1E�=Ev�D�$6 ���H� _FI+!�9�CORD� �_"36�r�B�1� �$ZDT�5�|"�%�4 *�L_NA�!(0�B:5DEF_I�H�B`6 TF5�96$962SF5@U`6IS��l��!���94ySF3T�]$4=��r"D �b�T,#�Dh�O��"LOCKE��C:?L?^7{QB@UME�BD2S D@UD�R&Bc%ES &DPT&B&{f{Q1C�  �1E�B1E2S1C�g�eH� P� iT� uQ���� W�X�e�S-���TE�a�$� }�LOMB_r�/w0�VIS��I�TY�A$�O�A�_FRIWs� SIuQYq��R%0�w00R�w3E#�W\xWh{Ț�^vn�_�y;AEAS�;B5�Vtŀ�P�2��v4~y5~y6�ORMULA_I����G�G� h �S.7e%COEFF_O1o r�1C��G���S�~"CA����/�#!GR�� � � $�P4F�"X� TM�W܄`�U2�S���#ER� qT�T�D�@�  ���LL<D�PS�_S�V�TH�$v�@��� G��@� ΂SwETUuSMEA�0��0��!�B�� g� q�] g �@����µ��Q���BH(0�Q�Q�T���qFB�f1�P�Q�P��t��� �0REC�A:���!SK_���� P�1_USER/�N�? s�N�/VEL�N�? �v�j��I�@� �M�T�!CFGD�� � *0� ONGORE�� ���� ~��� 4 ��8�XYZ�C��@ J#�ʠ_ERR��� ����!�0����2!:���� B?UFINDX�Ȣ��pR� H�CU��!_��1�A��<��A$Lt�AOQ咻�@ ��GĂ�� � $SI`;��p�0{R�VO��<���POBJE�����ADJU�"´ѰA�Y�AɳD��OU��@�_��1�B=�^�Ta .�v�-ǡ"DIR2�:�� ��ziGDYN�ry�v�T ���R^q� ����O�PWOR�� ��,� SYSBU���SOP��4�_���U�ˡ P�P���ŃPAQ������OP/@U����)"�f!�IMAG$���&�"IMw�@�I�N�p�?�RGOVCRDk���R��PЀ>�i� �`�S��L��PB�� ��PMC�_E�@4�[!N��M���f!_"1d"� k�S�L��E�� ��O�VSL�S�bDEX�QNP �2g ��_k��a@l��a@"�7�2�_"W�CZ�@�xf�4�l�_ZER��8�Ӄ�D�� @נ��3O�@RI±D
 ��0�����ǡ�ܰ�LD��Z�T A�TUS��u!C_TV�C��B����Ṕ��Se!���@E�� D �!���s�v3�A?�$���XE���\�p�;��㲠��U1PPoQPX�0.���]$3��7��P�G�����$SU�B��3]a����JMPWAIT��'��LOW�1���CCVF�1+0RK�,��&CCi�Rm�2�_IGNR_PL^��DBTB PsQFBW�0U��U� �TIG�j0IT'NLNS�R���R�]pNj0��PEED|��	�HADOW ��ʰE�����PSPDD�� L��A'�P"�0U!N���.��Rw�q�LY�@�  ���P4��D���$����f0� LE��� PA �P���xP�~}�S�ARSIZ�4�@�CMQܰO>@�9�ATT���-�����MEM�"f!�TU1X��}�qPL�0��� $���aSWI�TCH	�!WͰA�S��1"LLB�~�� $B�A+�D�S�BAMв�[Å)��w J5�����"6�&Y!_KGNOW��"k�U�#ADz(��-DQ��)?PAYLOA���`B3_D�7��7Z3�L]aA��>PLCL=_� !}�D2P�!��Q4��_6Fi9AC�?:��B4[�I?8!R�?70�[4B�p��Jq��1_JI1i���AND/�
��4I2�]1���qPLh AL_ �= -���!T��<pC�D3E���J3�0F� TU�PDCK��rR��CO��_ALPH CfCBE��(� O2L������� �s �� ?D_1:5224D��ARc��H��E�F�C��TIA4�Y5Y6�MOM�q�S:S'S:S4S��B% ADS^V'S^V4SPUB��R?T�U'S��U4R���@G@��/  �M,2�� �1!A��?� e$PIm����CZ�7i`�'9iI
kIkI+c�T�\f��\f����\Bg�W����HIGL#�& �f&\ K��f�c�h\�i\&SAMPk�d�t�gs&� �3 o�Fq�� z�Ut��_v�@ny�@ z�����P]u�q�b]uIN�|�p�c�x�{�t�&�z�x�t�{�GA�MM�uS
���$GGETW�@���D�D���
��IB���I.�$HI�_[�D�$z���E����A������LW��̆Ì��������B�f� AC�C�HKyг�ڐUNI_�`����B�H�q�u�Y�RS��|VX�GC ��$BH 1����I��RCH_D`X�����G��LEv��Z���嘩H���� M�SWFLV�QSCMR��10���SN�Wr3��:�|w�PnyxN�]�PI3A�VMETHO}モ�V��AX��h�X� ����ERI��t3�C�RB�5	�a�@FH4�q\s��ks���LĐq�OOP�\q��0�kq��APP��F�И4�U�@�&�sRTբ�O�0����a����T`1����T`஺+`��)�M�G��,&SV~��PD�G� ���GRyO� ��S_SA�!X��ū�NO�@C�� ��D�b��O?%?1h��o�W`�"_e���CDOA_�� UvP��u �h��g��h���æH3 >A0 M�U�o � ^�YLc�1�w��S�2Q��b�(����1��nӽ1�_đC�Z�M_W�A��� �w����M@j ��d0��A3)��	(����PM��R� � $Y�m��W"�n�԰L!51"� �D �D �D �4D{ ���N� d�C#���pXjO�C�qZ���P0 ��T� ���M�� W�T�f�xϊϜ�P���ّ�,#�A_��� |SA���:Yl�'Sl� 4S�Z����-ZR!\�P*!c!P���* 60�P�P��PMON�_QUp � =8�QCOU���`7QTH� HO[� 7HYS�ES�" �UE �xO5$ŋ  ? P �|�3�R_UN_TO��A�9O�b�P� P� `�C��/���INDE>��ROGRA��' �o�2��NE_NO��`IT�Q� D IwNFO��� ?!h�
�m��@�OI��� (p�SLEQ��f��e� ��D S�2��� 4�E�NABN�^ PTI�ON���ERVE�db[rac 3GCF.<� @ J�УqVh�h�R�\xn,"�PEDIT��'� �/��K�Q�c5��E��NU���AUT.��COPAY�Q�`,ra:�M���N +*�PRUT��R "N�OUC��a$Gep$��R�GADJ��� hS@X_��I͓���&���&W�(P�(�&�c� �N�0_CY�CN��QRGNSr8�P��`LGO7��s@NYQ_FRE�Q�RW�p�f-1SIZK8�LA��$1�!85S�p�eCREo���f8�IFa�NA q�%k4_G��ST�ATUS�VMA�ILrbA�1�L�AST�1aA�$EL;EM<� �9�FFEASII�Kr D�t��2���F٢�pn�I� l�$2�a��L�KBAB2�@E� r�`V�1cFBAS�B�dEn��QU�`�`'��${A�GRM�PR EC�qؐ�C���`��1��D.2�S�[�	~"B 2� �s ���tV�BW�B�Њp��ѡB3W�WߔDOU��ӔO��$Pݡ�@ОGRID�2B�ARS�gTYJ	��AOTO����� Q_�4!� �RnT�O��9� � ����POR��S��.�SSRV�0)�T�VDI0�T_e``#dPr`-g`-g4+i5+i�6+i7+i8a�F�?�<�O $VACLU~C�D@0}F8�� !E�;��S�1�۠A�Nõb�1y�12ATOTAL_�4I@r�PW3IvQ(tREGGEN&z;r��X�H`u����f��TR�C�2&q_S��w;pأAV�!��rsdBE�3�ݠB`��cV_�H�PDA��p�pS�_Y6���>6S�A�R��2� h"IG_SE�p�R�5�_d �tC_�V$C�MJ�C�T�DEE��b�I:�ZS�-�N1zC FB�HANCO� p�AG�2A3�qINT`�!��yFZ��MASKʣ�@OVR����ݠ���1��WV/ߠzT��A�_'Fd{�V�PS�LG%��a� \ ��?57��p�0S8���4f�Us�V�|��s��7aUP�TE|���@� (cq⟦J3�.�N3IL_�MM4�VQB۠��T!Q�𖣷�@C����5V�C-�P_�'��7�MN�V1M�V1�[�2j�2[�3j�3
[�4j�4[�����ޣ��ޣ����IN��V�IB�'�����2��2#�3�3#�4�4#���6�O�2����D`�Q`����P�L�0TOR ��I�NƵ��R��L���T $MC_F,  5���L ����pM?�I���OS� ]��f���KE�EP_HNADD" �!B�h@L�C�ᐐAbĮQ�t�c�O��A� ���pcë�c�REMz�bĺ1�R��Զ���U�4eb�HP�WD  B�S�BMӁ�PCOLL�AB���`e�qq2�� IT0��&"NO�FCALE����7� ,��FLK��A�$SYN��`�M���C@���pUP_�DLY���ODE�LA�л1�2Y��A�D����`QSK;IP$�� ��Pb aOp਒(���P_b  ��ד ��� �׵ � s �D`��Q`��^`��@k`��x`�څ`��9�!O�J2R� ���AX�@T'3���A���� >¡�>���RD�C�aT�� ��R�˸R`1ɺȲ
T�RGE�4CгXRFcLG���ŐSWX�
TSPC��!UM�_��ؓ2TH2N�RQk�� 1ݏ 	���Q8 � D� ��:�l@O2_PC�#��S��|�A.0L10_CL2�RC��́ � � b�'`����F(�� ����� ��+U��@г+� �b9�lC� �������~DESsIG��'UVL1���1��Hs10��_�DS�(����p  11�� l3�i���o�F&�AT��q$]Q07�'+$�  ��x����HOME�й2�������! �3��DVhz��� �4�������	// ��5��>/P/b/t/�/�/S ��!6��/`�/�/�/?? U
�!7��8?J?\?n?(�?�?38��?�? �?�?�?O-%S���  �A�Pp�6���E�T� aT���D	v�CIOՑ��IIp@5�OB�_O�P�ESr�C/!PO{WE��� �@�_п��"t �Z�BR$DSBf�G#NAOs��Cq�`�Q���Z�CIk _T_SPE%�z�CMD�W/ Â�a��ޘ�DBG_\@PU������SEq�̀ �2�4C=�'2S23�2�E� ���7E|o���ICEUSs<�U�ARIT�qq�OPB.ЭbFLOW�TR�@r���PƮaCUV` �aUX�Tҁ�a��ERFAiC;d��U�`�2wSCH��� t3�0���QH�@�$�p�pOM���A�  t���UPD����qPT�@Y�EX��x�c!�FA�e�G��r>fq � �цpZ�� (�AL� ��3u���:R;�  2�� �S���@��	� �$X���_�GROUQ�sT�\ ��vDSP�vJ/OGLI�cF����,a7�N�����ސ�f=K�`_MIR�q�Tf�MT��AP�`�c�*�Z�`�SYq��t�]��@�BRKH��avl�AXI~A  f�@�q��rρ�<�u�BSOC�v���N��DUMMY1�6,�$SV��D�EQnSFSPD_�OVR.����DL؂�sOR�P@N��b�Fv���pOV�u;SF�RUN����F8��a�sUFRAvN�TOldLCH�Ҍ���OVׄ8��pW�- ��sy�P�����_�8�� @E�TI�NVE$PKAOFS2ǐCSp��WD ���`�����R#�ÀTRO��R(�FD��(�M�B_C4��B� BL~���q0�6��qP�V�adB�` ���G1�D�AMB�$��`r�����_MH��b<��C���T$����q~CT�$HBK�a/�ءI�O_E�Q��PPA۪�������R��DVC_�PdCI�@q`RI�҆a`�1h���`�3h���"��`��pׁUdC�p�FCAB��^B[�"��&�k��h�O�UX/�SUOBCPU_R�pS�� ���Z��`��I�Z��?R��$HW_C@� t`���N��N@�pNp�$U-�z�|t�m�ATTRIEМ���pCYC��ұC�A���FLTR_2_FIqCsY��fVz��P�{CHK_�`�SCT�F_m�F1_w� ҉�FSeQR�r�CHA����A�Q�{b@�RSD��bQ��s`QP_To�? ��L�q`EM�@��Mn�T.��Np.��Ӷ��DIAGuRAI�LACV���MpL�O��f�<�$P�S�r`B �����P�RJ�SZ�& �Ct<�C 	��FUN��aRIN�Z�Y@0��?�pa��S_�pu àh�@Ѥh�-�Ѥ?CBLCUR}��aA������DAx�0i�����LD�`ˀ�����qr� ���T�I��}�Np$C�E_RIA��oRA�F�P�SG�[ L�T�2��Cs��C�OI<��DF_L�@P���as`LM�SF;H�RDYO�ѐRG� �Hb��Y@����MULSE����Ǽ�.s�$J�J�����FAN_ALM�MWRN!HACRD`@�ffs�2�Vaz�R�_��/�AU�R�R3ԇbTO_SBRU��p�
m�>�|G�MPINF���������REGF`FNV�`�Sb�DP�N�FL_Ž�$�M�����c��Np�(/C�P� ��b�h�PӐa��@$qAg$Y�R�a}r~�S�� �7�CEG�@�sˀ�A�P�D��25�����D�wAXE�wROB�z7RED�vWR�Pk�_���SYh��Ϡ:&S!'WRI�P�M�STOP�s�`l��%Eo��@�6��f"�pBa ��h&7�ӝ��OTO��@Y�ARY�s�"�ѝ��B�p�FIM��s$LI�NK��GTH�"�
pT_^#���8����!XYZ�b�*9�&OFFŐ�"�P� J�(� B�p4�D40��mP�`E3FI��^7�K�nSÄ4��t_J ,aNr���#��[ w$�*30��9`Е1���2�C#Q4�DU�³�3\%���TUR X"�E�!�X0 `�7FL� l�̳�$@5d)�35�Ғ 1�
�@K�pM/��6���p����cORQ�֠�qn�8��J�O N���E���q��DOV	E�AqM�`�Aj
U p
Uv	VaWαWpTANE��!
QL� r�A�IP��QU�A�W�Up�U.S�qER�qr�	 �E��Dp��TAQNpa5`��0�'��׶��AX��Nr �ᝰV��"+e��7i�� 7i��6j�6jq 6j�  6j� 6j06j1�06f ��3i��Ci��Si��ci ��si���i��i��i��i�a�iDEBUE�$@�L��tqڒ��"AB��ء ��CV͠D� 
�rq�r �u5��w���w���w� �wq!�w�!�w�!�w1�R��0L��"E3LAB�[2�EA�N�GROh���2E��B_�� �VM$��U0� l����E8��y��ANDr@ �@�T���%�Qy� ���M^ �������� NqT, ��+�VEL���eT5���=���E3NA�c�� �$��A�SS  ��i����� x��ʐSI����.��㆔�I���������AAVM, K� 2 ��� 0  �#5������%� %�	H�9�\������J���n��� 8�����G�������АBSQ� 1���� < �Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ��������������/�A�S�e��L�MA�X��Vh��5�  dz�IN����y�PRE_EXE��!����D�����А�IOCNV*B�� ȑ�P���0��1��wIO_�� 1ݛP $͠�r�]��Z��?�h���}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?��Q�c�z�LARMRECOV ������6LMDG �FQ k�LM?_IF F�� h��"�4�F�T���w���ϛϭϾ�, 
 ����b�n��1�C�T�$��x�_ߜ߀[����������s�NGTOL  ��� 	 A   �>�P�z�PPINFoO Ż Ķ�������   �»��者�����6�  �2�l�V���z�����������(: L^p������غPPLICAT�ION ?-������ArcTool � 
V9.1�0P/30O��?
88340-sF0S@105�-"47DF1x(�None��FRA� �6p�_ACT7IVEp�  �7��  �UTOM�OD ��5��CHGAPONL$/� 8#OUPLE�D 1�� �u y/�/�/�CUR�EQ 1	�  UT�)�,�,	�/�	5� 4���"_�ARC We=l��AW���"AWTOPKS6HKY?���/�/�/ ?v?�?�?�?�?�?�?  OOO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ�� ��(�:�L�^�p��� ܟ����ʟ�� �� $�6�H�Z�l�~�د�� ��Ư����� �2� D�V�h�z�Կ����¿ ����
��.�@�R� d�v��ϚϬϾ����ό�̹%TO(�/#DO_CLEANE/|�|�NM  -� �/������ ���.DSPDRY�R��V%HI" ��@ ��~������������� �2�D�V��MAX� c��1T't��Xc�sp"s�PL�UGGc d�p#%P�RC5�B�����m�_���O��>��SEGF< ^0.7 �߶�~������1LAP[�n03  2DVhz�������TOT�AL����USENU[ h+ I�M/2�� RGDISPM�MC^021C+3'�@@�"h$OY�{��I�RG_STR�ING 1
4+
_�M- S��
�!_ITEM1�&  n��/? ?%?7?I?[?m??�? �?�?�?�?�?�?O!O�3OEOI/O �SIGNAL�%�Tryout �mode�%In�p�@Simula�ted�!Out��LOVERR~X� = 100�"�In cycl��E�!Prog OAbor�C�!�D?status�D�@�cess Fau{lt\AlerT�	Heartbe�aSgCHand BrokeZEWOY_ k_}_�_�_�_�_�_�__��+_��/�_9o Ko]ooo�o�o�o�o�o �o�o�o#5GY8k}�_WOR: �+ �q)o�����%� 7�I�[�m���������Ǐُ����!�3�PO�+1QY��{B�|� ������ğ֟���� �0�B�T�f�x�����p����үT�DEV\� ��p��$�6�H�Z�l� ~�������ƿؿ����� �2�D�V�h�z�PALTm���{� ���������#�5�G� Y�k�}ߏߡ߳�����p������GRIy� �+E���m���� �����������!�3� E�W�i�{�������3�+ Rm��]���# 5GYk}��� ����1C<U��PREG�Ύ g�����/ !/3/E/W/i/{/�/�/��/�/�/�/�/[M�$�ARG_�pD ?�	���<1��  	�$[F	[P8]�P7�[Gq9/0SBN_CONFIGj@�<;�A�B�1�1C�II_SAVE � [D�1�3/0TC�ELLSETUP� <:%  O�ME_IO[M[L%?MOV_H�0	O�OREP��ZO%:U�TOBACK�1�<9�2FRA:\{ eO{�0�'`�@{�H�� �K�0 �23/08/13� 15:18:50{r8{_-_Z_Q_�L��z_�_�_�_�_�_�_{��_)o;o Mo_oqo�oo�o�o�o �o�o�o7I[ m�����p��!����  �A�_}C_\ATBCKCTL.TMH��`�r�������oKIN�I���E�5�1z@MESSAG�0ρ�1|D0ڋODE_D�0�6�5�O���wC�PAUSm� !��<; , 	��r0<5q��,		i�����ǟ��ß�� �!��-�W�A�{�e������D�N�TSK � T��O��z@UP3DT�͇d���XWZD_ENB8̈́�:'�STA̅<1��.1WJ@ODP�2�<;4W��)13-AU�G-2P7:33@P42O��˿ݿ�E{
{��߿*��7�`���o�03Dd� / a� �o�fϚ���j�ROoBGRPҨ�A��"�WEWEL�p���&id0�6-SEP����1�:0��E	LAB&��_2�{���9k�f��q�oߢ߯�������1C 57 ��f����ޭ�AXIS�0UN���Ԧ�1��� 	 ���Q��jE%�7z��_�~)Q�{V������D��1��t��{V����� �� -� ���� �?,������p����0�3�MET��2D鄰 PU�A�sQ�@��@��A�@mdA�A?����?&�>�E��=�i?I�6>��1?�@���5�SCRDCFG� 1<5�A ��5�2���@);M�O{Q�9 ��������^ �?Qcu��0 :'7}AGR=��X2��C�NA#@;;s	}D�_EDˀ�1�����%=-I�EDT-���m/����@!~BI/:�r2p_FB/�/  ���%2�/[/8?/��E�%??�/�/n?�/�#3�?6K�?O 7��+�?KO�?�?:O�?�#4�O�?�OO)N�O@_^OpO_�O�#5O_ �O�_�O)Nx_�_*_<_�_`_�#6o�_ho�_ )NDo�o�_o�o,o�#7�oWo4{o)N{ �o�oj�o�#8�'? ��*M�G���6���#9��̏ �h��)���Z�l�����!CR�/"���� X}r�ݟ$�6�̟Z��~% NO_DEL���GE_UNUS�E��IGALL�OW 1�� �  (*SY�STEM*L�	?$SERV_��L�~��POSREG���$£Lܗ�NUMxŪ�حPMUC�>L�LAYO�L��PMPAL|S��CYC10$��7�!�%�]�ULS�U�٭9� ��L�s���BOXORI�ɥCUR_��ح�PMCNV�晰10M���T4D�LIB����	*P�ROGRA��PG_MI%�O�a��AL/�n�X�a�B��ϗ�$FLUI_RESU=���ϯ�����MR������ ��Wr?�Q�c�u߇ߙ� �߽���������)� ;�M�_�q����� ��������%�7�I��[�6�LAL_OU�T ���#�W?D_ABOR>�g����ITR_RTN�  �Ā���N�ONSTO ��� O�CE_RIA3_Id���0 �� FCFG �*0��9_PA���GP 1CU������C;��� ��C�� C � (� M�C�8� @� H�  CUX� `� h� p� Ux��� �� �� �� �Rdv����?�HE�ON�FI����G_P6߰1C 1� ����/ /2/D/V/|h/�KPAUS��31��0 M�j/ �/���/�/�/�/?�/ 6?H?.?l?R?|?�?�?��?�?�?�?r,M��N�FO 1��}S  � 	�hOO;�=@B�7���yO  �'���Dd�8C���6���X �hB�@�d�����XD̿7�3���W���k3�gO=C��Ǹ�COLLEC+T_=+F��R�GEN/����R�A�NDE�C�G�R��1234567890[W:ұ�0SY_kV��
 %}�;�)�_�_���_�_o ���_�_Too1oCo�o goyo�o�o�o�o�o, �o	t?Qc� �������L���5V��2�K �]9RIO !DYQ����Ώ���l���TRr 2"��� ��
-����#��<��Y_MO5Rz�$w ��ŕ <Ařݟ˟��%�����m{�%��,�?$���x�;�K��;��� R=&�O����~��C4  A�����;�=A{�Czg  B�$B�"o  @Ң���;�:dڍ��ARIJ=S'��?�z�(����/�d��T_DE-Fz� X�%J�������NUS<��0���KEY_TBL�  �06B�	
��� !"�#$%&'()*�+,-./dW:;�<=>?@ABC�e�GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����h����͓��������������������������������������������������?������}!b��LCK��	b���S�TA����_AUT/O_DO��&��INDT��_T10�"�T2o��V� TRLd�LE�TE����_SCREEN ��kcscU� MMENU 1)�� <o�|�D� UE#�M��i�k��� ����������6��� l�C�U���y������� ���� ��	V-? e�u����
 ��R);�_ q����/�� <//%/r/I/[/�/�/ �/�/�/�/�/&?�/? 5?n?E?W?�?{?�?�? �?�?�?"O�?OXO/O AO�OeOwO�O�O�O�O�_�O�OB__�_M�ANUAL���D�Bc�j�����DBG�_ERRLj�*�D� Q_�_�_�n�QNUMLI�M��[���
�QP�XWORK 1+��__oqo�o�o�o�S�DBTB_�� �,�]ģ4����o�DB_AWAYz�SD�GCP ���=��1b�b_AL`��b�RY���ը���X_�P 1-��h�
No���|��f�_ML�IS�
{@|{��sONTIM�כ�����vGy
���\sMOTNEN�D��[tRECOR�D 13� �<���G�O���u� ��
r��ŏ׏鏀�� ���<���`�r���� 1���)�ޟM���&� 8�ӟ\�˟����� ȯگI���m�"���F� X�j�|�믠��Ŀ3� ����ύ�Bϱ�M� տ�ϜϮ���/���S� ��w�,�>�P�b��φ� q�߼�+������s� (���^��߂��� =����K� �o�$�6� H�����~������� �������� ��D���hz���bTO�LERENCtB��QrpL�͈PC�SS_CNSTC�Y 24?i��P�Or�	);Q _q������ �//)/7/I/[/��DEVICE 25� �f�/�/ �/�/�/??,?>?P?�b?��HNDGDg 6��`Czu:|O��LS 27�-t?�?�?OO,O>O�POv?�PARAM 8hy8rwUbD�5��5SLAVE �9�=�7_CFG �:�ObCdM�C:\� L%04�d.CSVaO"�c�	_!�>A 6SCH>P�1�bNI_~_�G�bFnR�Q�_�Y�Q�@JP��S�^"���a�>_CRC_?OUT ;�-�a~fO_NOCOD�@�<hw�MSGN �=^�G�#M��06-SEP�-23 13:0�19P�A13-�AUG~b5:19�9P�& Wz�z�i�abN�`ra�M���Þ�j���a�n�CVERS�ION ej�V4.2.11��{EFLOGIC� 1>� 	��X�@Iy�QY}+rPROG_ENB<�\�6ysULS�w �6�+r_ACCLI�M�v��C���sWRSTJNT0�F��A+qMO�|�Q�Pb�tINIT �?�
^��A �vO;PT�@ ?	6���
 	R57Y5bCc�74h�6i��7i�50��t��2�i��X��%wF�TO C R��o�&vV��DEX�wd�riP�$�PATH AejA\�q�����HCP_CLNT�ID ?	v�C ��[Zß�IA�G_GRP 2D��I > �	 @K�@�G�?���?l��>� �@ٚ��8�ٜ5��� |a�O�?�b�?> ���i�^?�Vm�?Sݘٙf�403 6789?012345������ �s���@nȴ@i�#�@d�/@_�w�@Z~�@U/�@O�@I��@D(�ٚѠiQ@Š6Tp6P�� A�� � 9PB4ٜP� ٔR�iQ
Т1���-@)hs@�$��@ bN@���@ڠ���@�D@+2�	��-�2�A�2��P�R��@N�@I�@D��@>�y@9���@4��.v�@(?��@"�\����𬿾�пV�L�@�Gl�@BJ@�<z�@6ڠ0��`@*�$����@��&�8��J�\�V�=q@���F@|��@33@�R�@-?����?��`?�+ �ϲ��������̑҂���-@&�@�����!?�?� �,� >�P�b�t�V� �(�:� �^�p���D���� ����x����6�H�&� l�~����:���q� ����ѡ�x�������Y���?�zy���(�5AF�4� ��L4�R� (�@�p�.8�Q�@-: I f�m@���%�Ah.��=H�9=Ƨ�=�^5=�v ��>�(�=��,��,�^� �iQC)�<(�U�R 4���[��ٙA@hR?0� ��"��0Vh4�� t�8����
/޴�>��y,"��R=���=��yz<!(���G�T/G�(�8U8U����($@9P��*���uB�J���B��B��B%�!(��T�/�.'�p5�.�*11n,�\@��=�-��c+�a Bk �B��BC�A��@�pZ?؟�?iQ<�P�  3>��?y?O��3P�1��3\�N�2�Jd��0�18���BDd�8C�3Qu��?O OD9O�(TOZBٙ�9�6���.�B� R�)O�O�O�O�O�O�O|__>�{Dٙ>�� ����'_u_�CT_CONFIG EDo>�ceg�U��STBF_TTS�w
�y�S p�s��V5`MAU�p��r�MSW_CF�PF���  )��jOCV7IEW�PG'm3���ןyo�o�o�o�o �oPrgo�o 2D V�oz����� c�
��.�@�R�d� ���������Џ�q� ��*�<�N�`�� ������̟ޟ��� &�8�J�\�n�������`��ȯگ�|\RC c	H`��R!����$�Y��H�}�l�����ſdS�BL_FAULT� I�<h߱GP�MSK�W�PTD?IAG J�Y�!��S��QU�D1: 6789?012345O¬RC��W��Pb_�ϝϯ� ��������	��-�?� Q�c�u߇ߙ߫�j�?����
z��߂VTR'ECP(�:�
H�:� a���y�v����� ��������*�<�N� `�r��������������=gUMP_OPT�ION�P���TR� b�S�PME��UY_TEMP�  È�3B�Q0m �L1WUN�I`�Um�YN_?BRK KRo=f?EDITOR���F�_�ENT �1L�  ,�&	LABWEL�D_2����&M�AIN @&
� _�5fM20���ֲ��� �/�/C/*/g/N/ �/�/�/�/�/�/�/�/ ????&?8?u?\?�? �?�?�?�?�?�?O)O�OMO4I� MGDI_STA�+am��NCsC1M'k �����O�O��
��d ��_'_9_K_]_o_�_ �_�_�_�_�_�_�_o #o5oGoYoko}o�o& �o�o�o�o�iQ�o "4FXj|�� �������0� B�T�f�x��j�o���� ͏ߏ�o��'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uϏ�}ϫ� ���������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m�ϙϣ����}��� ���!�3�E�W�i�{� �������������� /ASe�� ������+ =Oas���� ���//'/9/K/ ]/o/��/�/�/�/� �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgO�/�O �O�O�O�/�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oyOko�o�o�o�O �O�o%7I[ m������ ��!�3�E�W�qo�o ������Ï�o���� �/�A�S�e�w����� ����џ�����+� =�O�ɏ{��������� Տ߯���'�9�K� ]�o���������ɿۿ ����#�5�G�Y�s� }Ϗϡϳ�ͯ������ ��1�C�U�g�yߋ� �߯���������	�� -�?�Q�k�Y���� �ϻ�������)�;� M�_�q����������� ����%7Ic� u���Y���� �!3EWi{ �������/ ///A/[mw/�/�/ �/��/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO e/oO�O�O�O�/�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCo]Ogoyo�o �o�O�o�o�o�o	 -?Qcu��� ������)�;� UoG�q������o�oˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�M�_�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� ��W�a�sυϗϱ��� ��������'�9�K� ]�o߁ߓߥ߷����� �����#�5�O�Y�k� }��ϳ��������� ��1�C�U�g�y��� ������������	 -G�5cu��� ����); M_q����� ��//%/?Q[/ m//5/��/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O7/I/SOeOwO�O�/ �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'oAOKo ]ooo�o�O�o�o�o�o �o�o#5GYk }������� ��9oC�U�g�y��o ������ӏ���	�� -�?�Q�c�u������� ��ϟ����1�#� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���)�;�E�W�i�{� ���ϱ���������� �/�A�S�e�w߉ߛ� �߿���������3� =�O�a�s�ϗ��� ��������'�9�K� ]�o������������� ����+�5GYk �������� 1CUgy� ������	/# /?/Q/c/}s/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�?��?�?O/ �$E�NETMODE �1N~%��  + + �&%HOZK*@RROR�_PROG %�7J%%&�O�IxETA�BLE  7K��/�O�O_WxBSE�V_NUM FB?  �AA=P�xA_AUTO_ENB  dE?CuDw_NORQ O7K�YA<R  *�*�P��P��P��PHP�+�P�_�_�_nTFLsTRZ_lVHIS9S�)!?@g[_ALM �1P7K �&$�\% +�_no�o�o��o�o�o�__2RtP  7K�QZBz*@�TCP_VER �!7J!�O�o$E�XTLOG_RE�Qf�eY_sSI�ZhZtSTK�y��U�\rTOL � )!Dzb�{A Zt_BWD�``�p�V�q_B�sDI�qw Q~%�sxXD)!�{STEP���*@0�OP_DO��(AFDR_GR�P 1R7I�Qd �	��Z@��n&����c?���$,MT�� ��$ ����ن�������B����CF��C ���CP�Bԟ�B��H`�A��0�A��B��]�B)�jA�WA���� ��r�]���������ޟ�ɟ  @�?�A���>(��A��`�
 K��uA�	�)!A��r�Eb؟ҟw�b�䛯*�@7���@�3�3@�Ǡˣ�@�¡毄�����F;@ 5�E��@�5��%��L�FZ!�D�`�D�� �BT��@��Þ�?�  ��#�6������5�Zf5�ES�������E�K$F�EATURE �S~%�p^A�ArcTool ��)"Engl�ish Dict�ionary*�4�D Standa�rd#�Analo_g I/O"�A5�e Shiftw��rc EQ Pr�ogram Se�lect��Sof�tpar�ǝ�We�ld��cedur�es���Core����Rampin�g_�uto��wa~�Update(��matic Ba�ckup(�V�gr�ound Edi�t �-�Camer�ar�Fv�Cell�r�{�nrRndI�m[Ӓ�ommon� calib UI����sh������1c�	���ne�	�Kty��s����nt����Monitor�=�ntr�eli�ab��)�DHCP�˒�ata Ac�quish��ia�gnosR�o���o�cument V�iewet��ua���heck Sa�fety��-�ha�n�� Rob��r�v��q!���)�F�s���F���-�xt oweavS�ch%�xt. DIO���nfi"�|�end..�Errs�L���Ji�s��rm��� �p�'�FCTN Me�nu�����TP ;In��fac�-��Gen��l��Eqs L��8igE'�9m�p Mask� Exc*�gr�H�T% ��xy Sv���igh-Spe.�Ski�ԍ��~��mmunicQ�{on��Hour ����s�(conn�X�2�ncr' sGtru>��
!e����J��-�KARE�L Cmd. L� ua�XRunw-Tiq�EnvN���:�+U�sS�S/�W*�Licens�e�����Book�(System)�'�MACROs,~�/OffseZ��MMRm�i���Me�chStop��t������i���1&x�.�o�S�D.od��wCit��g(i���.���+Optm�/#��'fil��'g��?ulti-T  ��+�ORNTBAS�E Fun+-�P�CM f"8(�Po���� �I=Regi2�r��,6ri��!9~9p�Nu����8��Adju� �>���=tatu}1�?��n,�RDM0�ot;��scoveD�)Ee�a� q�Freq �Anly��Rem' ��nR�)E5B5�N9�ues�ńGo���r )�SNPX b�#�SN% Cli���N��P rC��OU�Q 8$P�Eo�t ssag յE����O!p 0��V^/I|&]UMILIB�_~`RP Firm9�:p^PAccn�v��TPTX��^Tel�n��_aQ��q]o�r�@ SimulQar��!fu��P8��XZmЍ�#&��ev�.]U1�ri��_?USB po�����iP��a��fR �EVNT�o�`nexcept.�j@W4X�ej�P�VC��r��-(V��.r�_?u�K�9{S�@SC�UqS�GE�|uUI&�Wx��8�|b PlF �~5���� (���������6�uZDT Appl�'��f��s�Grid9AplCaym�mPZԇ�R%r.R�����F� A��200i��c�la�rm Cause�/h@edE�Asc{ii��Load���1�UplG���yc���~�0�`� RA�e`���yQ�NRTL��_4nline Hel��-6',6{0�x1��tr"�64M?B DRAM����FRO �����c� tPB� .'�mai����K�RR�6L��Sup�b�!}9à��} croL4C�E��9v#rt�4C&���z� .�@�m�d�v������� ٿп����3�*�<� i�`�rϟϖϨ����� �����/�&�8�e�\� nߛߒߤ��������� ��+�"�4�a�X�j�� �������������'� �0�]�T�f������� ����������#, YPb����� ���(UL ^������� �//$/Q/H/Z/�/ ~/�/�/�/�/�/�/? ? ?M?D?V?�?z?�? �?�?�?�?�?O
OO IO@OROOvO�O�O�O �O�O�O___E_<_ N_{_r_�_�_�_�_�_ �_oooAo8oJowo no�o�o�o�o�o�o �o=4Fsj| �������� 9�0�B�o�f�x����� ��ȏҏ�����5�,� >�k�b�t�������ğ Ο����1�(�:�g� ^�p���������ʯ�� � �-�$�6�c�Z�l� ��������ƿ���� )� �2�_�V�hϕό� �ϸ���������%�� .�[�R�dߑ߈ߚߴ� ��������!��*�W� N�`�������� ������&�S�J�\� ���������������� "OFX�| ������ KBT�x�� ����///G/ >/P/}/t/�/�/�/�/ �/�/???C?:?L? y?p?�?�?�?�?�?�? 	O OO?O6OHOuOlO ~O�O�O�O�O�O_�O _;_2_D_q_h_z_�_ �_�_�_�_o�_
o7o .o@omodovo�o�o�o �o�o�o�o3*< i`r����� ���/�&�8�e�\� n���������ȏ��� ��+�"�4�a�X�j��� ������ğ����'� �0�]�T�f������� ��������#��,� Y�P�b�|��������� �����(�U�L� ^�xςϯϦϸ����� ����$�Q�H�Z�t� ~߫ߢߴ�������� � �M�D�V�p�z�� ����������
�� I�@�R�l�v������� ������E< Nhr����� �A8Jd n������/ �/=/4/F/`/j/�/ �/�/�/�/�/?�/? 9?0?B?\?f?�?�?�?��?�?�?�?�1  H541�3zA2FR782 G{50 EJ614DG{76 EAWSP,G]1[GRCRPH8\F{TUgFJ545DH�[FVCAM ECL�IO�FRI�GUI�F,F6�GCMSC��HgFSTYLDG2ދFCNRE,F52�[FR63+GSCH� EDOCVLVCS�U EORSFR8k69DG0OG88FwEIO�FR547F�R69[FESETt�GrGJqIWMG�GޒWMASK EPRkXYX7 FOC�FB�P3�H7F�PCH3f[J6BH53{VHEhwLCH�VOPL�V�J50/fPS�gM�CfG�`�W55OFMgDSW�g"gOP"gGMPR�F<PSh0CFoORBS fCM�G�0w�POG50Sg5�1�G51Ox0�FP�RS�W69fFR�D�FFREQ,FMsCNVmXH93CF�SNBA�GFgSH�LBVM�w<P3WNuN_h2CFHTCgF�TMIV4@{VTP�A�FTPTX(�EL�v�`{W86G4@FwJ95�FTUT#g�95fUEV�VU�EC�VUFR�FV�CCψOFVIP�VCSCW�CSG�'VaPI�hOFWEB�gFHTTgG62WWkIO�Ry�CG:��IG�IPGvI�RCVDG"gH7]5�FR66��7�WURMz2/fR]j4fp��OF�@FNVD�V�D0��F�ALOn�VCTO�GNNf�M}xOLXEND:,FLڇFVR�E�8 ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿���  H�541��2#�R�782$�50$�J�614T�76$�A�WSP4�1s�RC�Rd�8t�TU��J�545T�s�VCA�M$�CLIO��R]I��UIF4�6���CMSC4܃�ST�YLT�2��CNR�E4�52s�R63�3�SCH$�DOC�V��CSU$�OR�S��R869T�0vc�88#�EIOC�wR54C�R69s�OESET�˒�J���WMG$��MAS�K$�PRXYd�7&$�OC�`�3��Cʴ`�S�3��J6R�5u3��H�LCH��wOPL��J50��PSb�MC��p�c�{55c�MDSW��v��OP��MPR�����0S�ORBS��CM#�0`�c��50�51��51�c0��PRSS�6�9��FRD��FR;EQ4�MCNT����H93S�SNBA�$��SHLBT�MX2�Г�NN#�2S�wHTC��TMIc��@���TPAC�TPTX�EL�
p���q8B�@�#�J95�ʷTUT��95��U�EVS�UEC��U�FR��VCCc,O��VIPc�CSCN�CSG����Id��c�WEB��HTT���6��WIO�*R��CG�+IG�+I�PG#
IRCc�D�G��H75��R6U6�;7B�Ra2��R!�4��0c�0�#ʷNVDS�D0�;F�!LALO��CTO���NN��M�OL�R�END4�Lr+FVRC�ȺO�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o �o�o�o�o�o0 BTfx���� �����,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������0 BTfx���� ���,>P bt������ �//(/:/L/^/p/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� �}�STD�?LANG(�#� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������ +=Oas��� ����'9�K]o��RBT'�OPTN���8��
+DPN&�"/ 4/F/X/j/|/���/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z?  ��?�?�?�?�?��?�=99E�$�FEAT_ADD ?	���/A�7@  	 �8@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n������������������""DDEMO� S/I   �8i_q�� ����
- 7d[m���� ��/�/)/3/`/ W/i/�/�/�/�/�/�/ ?�/?%?/?\?S?e? �?�?�?�?�?�?�?�? O!O+OXOOOaO�O�O �O�O�O�O�O�O__ '_T_K_]_�_�_�_�_ �_�_�_�_�_o#oPo GoYo�o}o�o�o�o�o �o�o�oLCU �y������ ���H�?�Q�~�u� ������������ �D�;�M�z�q����� �����ݟ�	��@� 7�I�v�m�������� �ٯ���<�3�E� r�i�{�������޿տ ���8�/�A�n�e� wϤϛϭ��������� �4�+�=�j�a�sߠ� �ߩ����������0� '�9�f�]�o���� ����������,�#�5� b�Y�k����������� ������(1^U g������� �$-ZQc� ������� / /)/V/M/_/�/�/�/ �/�/�/�/�/??%? R?I?[?�??�?�?�? �?�?�?OO!ONOEO WO�O{O�O�O�O�O�O �O___J_A_S_�_ w_�_�_�_�_�_�_o ooFo=oOo|oso�o �o�o�o�o�o B9Kxo��� ������>�5� G�t�k�}�������͏ ׏����:�1�C�p� g�y�������ɟӟ � ��	�6�-�?�l�c�u� ������ůϯ���� 2�)�;�h�_�q����� ����˿����.�%� 7�d�[�mϚϑϣϽ� ��������*�!�3�`� W�iߖߍߟ߹����� ����&��/�\�S�e� ������������ "��+�X�O�a����� ������������ 'TK]���� ����#P GY�}���� ��///L/C/U/ �/y/�/�/�/�/�/�/ ?	??H???Q?~?u? �?�?�?�?�?�?OO ODO;OMOzOqO�O�O �O�O�O�O
___@_ 7_I_v_m__�_�_�_ �_�_o�_o<o3oEo roio{o�o�o�o�o�o �o8/Ane w������� �4�+�=�j�a�s��� ��ď��͏����0� '�9�f�]�o������� ��ɟ�����,�#�5� b�Y�k���������ů ����(��1�^�U� g������������� ��$��-�Z�Q�c�}� �ϴϫϽ������� � �)�V�M�_�y߃߰� �߹���������%� R�I�[�u����� ��������!�N�E� W�q�{����������� ��JASm w������ F=Ois� �����/// B/9/K/e/o/�/�/�/ �/�/�/?�/?>?5? G?a?k?�?�?�?�?�? �?O�?O:O1OCO]O gO�O�O�O�O�O�O _ �O	_6_-_?_Y_c_�_ �_�_�_�_�_�_�_o 2o)o;oUo_o�o�o�o �o�o�o�o�o.% 7Q[���������*�!�M�  D�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������'|9K	  L Qgy����� ��	-?Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{��������� ������/APU Hk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A��S��$FEAT_�DEMOIN  �X�����X��k�INDEXx�����k�ILECO�MP T�������f����SETUP2 �U��Â� � N �_AP2BCK 1V��?  �)T�"�"1�%�U�X���C� ��V����;�П_�ݟ ���*���N�`�� �����I�ޯm��� ��8�ǯ\��i���!� ��E�ڿ�{�ϟ�4� F�տj����Ϡ�/��� S���w���߭�B��� f�x�ߜ�+�����a� �߅��,��P���t� ���9���]���� ��(���L�^����� ����G���k� �� 6��Z��~�� C��y�2D �h����Q �u
//�@/�d/ v//�/)/�/�/_/�/��/?�/%?N?ȉ��P� � 2�*.cVRU?�?0*�?��?
3�?�?�%�0PC��?#O0FR6:DOON�?sOKT�� �O�O8E�O�Lz�dO�O�&*.F�?*_1	:C_W\�O{_
[STM�_�_7B=@�_"�]j_�_
[H�_2o��W o�_�_�oZGIF�o�o�U�oaosoZJPG<�U(0�o�o�JJS���0Rs�j%
J�avaScript�CS�C��V�0�� %Cas�cading S�tyle She�etso�� 
AR�GNAME.DT��<�P\��p��q��󏟏�DISP*��.ބ9����	�i�w�#�
TPEINS.XML���Ώ:\��x�ځCu�stom Too�lbar��*�PA?SSWORDn��.?FRS:\>����_�Passwor�d Config ��/ȯW�����4?"� ��F�X��|������ A�ֿe�������0Ͽ� T��Mϊ�Ϯ�=��� ��s�ߗ�,�>���b� �φ��'߼�K���o� ����:���^�p��� ��#����Y���}�� ���H���l���e��� 1���U������� �� DV��z	�-? �c���.�R �v��;�� q/�*/��`/� �//}/�/I/�/m/? ?�/8?�/\?n?�/�? !?�?E?W?�?{?O�? 	OFO�?jO�?�O�O/O �OSO�O�O�O_�OB_ �O�Ox__�_+_�_�_ a_�_�_o,o�_Po�_ to�oo�o9o�o]ooo �o(�o!^�o� ��G�k �� �6��Z������ ��C����y����2� D�ӏh�������-� Q��u������@�ϟ 9�v����)���Я_� �����*���N�ݯr� ����7�̿[�ſ� ��&ϵ�J�\�뿀�� �϶�E���i��ύϟ��4���$FILE�_DGBCK 1�V��!���� < ��)
SUMMAR�Y.DG>���M�D:r߲���D�iag Summ�ary����
CONSLOG�ߋߝ����6���Console log7����	TPACCN�,��%y����T�P Accoun�tinX���FR�6:IPKDMPO.ZIP����
��;�����Excep�tion?����MEMCHECK�������J�Mem�ory Data����"l�)	FTP)������L�mment �TBDG�L >�I)ETHERNET<�΁�����Ethern�et N�figu�ra^���1DCSVRF;!3L���% verify allO��M.cDI�FFD*<���{%fdiff�����CHG01 ���V/a�~/�- )2L/3/E/�/�{/�/"3�/�/�/�^? �/�?6�VTRNDIAG.LS�?;?M?�?���1 Ope� �Log ��nos�tic���)�VDEV�2DA�T�?�?�?�?bV�isADevic9eOKIMG�21��AOSO�O�#~DImsag�OKUP/@�ES.O�OFRS�:\._o]��Up�dates Li�sto_���@FL?EXEVEN��O��O�_a�Q UI�F Evb	@�_ � ,�t)
P�SRBWLD.C	Mo��ZR6oq_K��PS_ROBOW�ELh�:GIG�E	Oo�_�o��G�igEXo�N��A�)�aHAD�OW�o�o�o|���Shadow C?hanges���a�<rRCMERRtYk �����pCFG Er�ror�@tail>� MA����pSGLIB���8��rI� St� A�-�>��)r�Z�D�o��o����Z�D@ad��3� <rNOTI��������Notif�ic�3�(f�AG ��������;��� _����$���H�ݯ �~����7�I�دm� ���� ���ǿV��z� �!ϰ�E�Կi�{�
� ��.�����d��ψ�� ��*�S���w�ߛ߭� <���`�����+�� O�a��߅���8�� ��n����'�9���]� �����"���F����� |���5��Bk�� ���T�x �C�gy� ,�P���/� ?/Q/�u//�/�/:/ �/^/�/?�/)?�/M? �/Z?�??�?6?�?�? l?O�?%O7O�?[O�? O�O O�ODO�OhO�O _�O3_�OW_i_�O�_ _�_�_R_�_v_oo �_Ao�_eo�_ro�o*o �oNo�o�o�o�o= O�os��8� \���'��K�� o������4�ɏۏj� ����#�5�ďY��}� �����B�ןf���� ��1���U�g������ ����P��t�	���� ?�ίc�򯇿��(��� L��󿂿Ϧ�;�M���$FILE_F�RSPRT  ���1�����\�MDON�LY 1Vp�(�� 
 �)M�D:_VDAEX?TP.ZZZN��������6%N�O Back f�ile ��(�S�6)ܿ7���[�$�h� ��ֿ��D�����z�� ��3�E���i��ߍ�� .���R���v������ A���e�w����*��� ��`�����+��O ��s��8�\ ��'�K]�����`�VIS�BCK��x���*�.VD�/pF�R:\�ION\�DATA\���pVision VD�./<v/�/ ��/��/_/�/?�/ *?�/N?`?�/�??�? 7?I?�?m?OO�?8O �?\O�?mO�O!O�OEO �O�O{O_�O4_�O�O j_�O�_�_[_�_S_�_ w_�_o�_Bo�_foxo o�o+o�oOoao�oV��LUI_CONF�IG Wp�|�{ $ �c��{p�Xj|����y@p|x�o�� � �2�B��e�w��� ����D�������� +�O�a�s������� @�͟ߟ���'��� K�]�o�������<�ɯ ۯ����#���G�Y� k�}�����8�ſ׿� ���϶�C�U�g�y� �ϝ�4���������	� ���?�Q�c�u߇�� �߽���������)� ;�M�_�q����� ���������%�7�I� [�m����������� ������!3EWi {������ �/ASe�v �����z// +/=/O/a/��/�/�/ �/�/�/v/??'?9? K?]?�/�?�?�?�?�? �?r?�?O#O5OGOYO �?}O�O�O�O�O�OnO �O__1_C_U_�Oy_ �_�_�_�_X_�_�_	o o-o?o�_couo�o�o �o�oTo�o�o) ;�o_q���� P����%�7�� [�m��������L�ُ ����!�3�ƏW�i��{�������A�͐x���ʓ�$FLUI�_DATA X�������D��RESU_LT 2Y��#�� �T�/�wizard/g�uided/st�eps/ExpertٟZ�l�~��������Ưد�������Continu�e with G7�ance�W�i� {�������ÿտ���,�� ˒-̑��><�0 �M�<������\��.�ps ϧϹ��������� %�7�I�[�m�,�M��� �߸������� ��$� 6�H�Z�l�~�\�N�`��r���torch ������*�<�N�`� r���������y����� &8J\n� ����������>��wproc��H Zl~����� ��/��2/D/V/h/ z/�/�/�/�/�/�/�/�
??��7?{����@�TimeUS/DST&?�?�?�? �?�?OO,O>OPObO~%�EnablE� �O�O�O�O�O�O__�&_8_J_\_n_˒�8�F?�_j?|?�624 �?�_o"o4oFoXojo |o�o�o�oqO�O�o�o 0BTfx� ���_�_�_�_w��-�?�Region �R�d�v����������Џ���!�America<@�R� d�v���������П����!��qy��P�8�$��2Edi��� ����ʯܯ� ��$��6�H�Z�+ Tou�ch Panel� �� (reco/mmen��)h��� ��ѿ�����+�=�O�a� ��0�B���f�|x��2acces/� ����/�A�S�e�w���ߛ߭�,Con�nect to Network�� ����)�;�M�_�q����$���p��ϚϬ��\!�ϐ0I�ntroduct >�Q�c�u��������� ������ /);M _q������� 0?��0 
��R#����� ��//(/:/L/^/ �/�/�/�/�/�/�/� ??$?6?H?Z?�x3P:H�?l�? �?�?OO+O=OOOaO sO�O�O�Oh/�O�O�O __'_9_K_]_o_�_ �_�_�_v?�?�?�_�? #o5oGoYoko}o�o�o �o�o�o�o�o�O1 CUgy���� ���	��_*��_N� ou���������Ϗ� ���)�;�M�_�p� ��������˟ݟ�� �%�7�I�[��|�>� ��b�ǯٯ����!� 3�E�W�i�{������� p�տ�����/�A� S�e�wωϛϭ�l��� ���ϴ���+�=�O�a� s߅ߗߩ߻������� �¿'�9�K�]�o�� �������������  ���D�V��}����� ����������1 CU�y���� ���	-?Q �Z�4�~�j��� �//)/;/M/_/q/ �/�/�/f�/�/�/? ?%?7?I?[?m??�? �?b���?�?�!O 3OEOWOiO{O�O�O�O �O�O�O�O�/_/_A_ S_e_w_�_�_�_�_�_ �_�_�?�?�?�?LoO so�o�o�o�o�o�o�o '9K
_o� �������� #�5�G�Y�o*o<o�� `oŏ׏�����1� C�U�g�y�����\�� ӟ���	��-�?�Q� c�u�������j�|��� 𯲏�)�;�M�_�q� ��������˿ݿ￮�  �%�7�I�[�m�ϑ� �ϵ��������ϼ�� �B��i�{ߍߟ߱� ����������/�A� S�d�w������� ������+�=�O�� p�2ߔ�V߻������� '9K]o� ��d����� #5GYk}�� `��������/1/ C/U/g/y/�/�/�/�/ �/�/�/�?-???Q? c?u?�?�?�?�?�?�? �?�O�8OJO?qO �O�O�O�O�O�O�O_ _%_7_I_?m__�_ �_�_�_�_�_�_o!o 3oEoONO(Oro�o^O �o�o�o�o/A Sew��Z_�� ����+�=�O�a� s�����Vo�ozoď� �o�'�9�K�]�o��� ������ɟ۟ퟬ� #�5�G�Y�k�}����� ��ůׯ鯨���̏ޏ @��g�y��������� ӿ���	��-�?��� c�uχϙϫϽ����� ����)�;�M��� 0���T���������� �%�7�I�[�m��� Pϵ����������!� 3�E�W�i�{�����^� p߂�����/A Sew����� ����+=Oa s������� ��/��6/��]/o/�/ �/�/�/�/�/�/�/? #?5?G?X/k?}?�?�? �?�?�?�?�?OO1O CO/dO&/�OJ/�O�O �O�O�O	__-_?_Q_ c_u_�_�_X?�_�_�_ �_oo)o;oMo_oqo �o�oTO�oxO�o�O�o %7I[m� ������_�!� 3�E�W�i�{������� ÏՏ珦o��o,�>� �e�w���������џ �����+�=��a� s���������ͯ߯� ��'�9���B��f� ��R���ɿۿ���� #�5�G�Y�k�}Ϗ�N� ������������1� C�U�g�yߋ�J���n� ���ߤ�	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������߮� ����4��[m� ������! 3��Wi{��� ����////A/  $�/H�/�/�/ �/�/??+?=?O?a? s?�?D�?�?�?�?�? OO'O9OKO]OoO�O �OR/d/v/�O�/�O_ #_5_G_Y_k_}_�_�_ �_�_�_�?�_oo1o CoUogoyo�o�o�o�o �o�o�O�O*�OQ cu������ ���)�;�L_�q� ��������ˏݏ�� �%�7��oX�|�> ����ǟٟ����!� 3�E�W�i�{���L��� ïկ�����/�A� S�e�w���H���l�ο ������+�=�O�a� sυϗϩϻ����Ϟ� ��'�9�K�]�o߁� �ߥ߷����ߚ��߾�  �2���Y�k�}��� ������������1� ��U�g�y��������� ������	-��6� �Z�F���� �);M_q �B������/ /%/7/I/[/m//> �b�/�/��/?!? 3?E?W?i?{?�?�?�? �?�?��?OO/OAO SOeOwO�O�O�O�O�O �/�/�/�/(_�/O_a_ s_�_�_�_�_�_�_�_ oo'o�?Ko]ooo�o �o�o�o�o�o�o�o #5�O__z<_� �������1� C�U�g�y�8o������ ӏ���	��-�?�Q� c�u���FXj̟� ���)�;�M�_�q� ��������˯��ܯ� �%�7�I�[�m���� ����ǿٿ������� ��E�W�i�{ύϟϱ� ����������/�@� S�e�w߉ߛ߭߿��� ������+��L�� p�2ϗ��������� ��'�9�K�]�o��� @ߥ����������� #5GYk}<� `�����1 CUgy���� ����	//-/?/Q/ c/u/�/�/�/�/�/� �/�?&?�M?_?q? �?�?�?�?�?�?�?O O%O�IO[OmOO�O �O�O�O�O�O�O_!_ �/*??N_x_:?�_�_ �_�_�_�_oo/oAo Soeowo6O�o�o�o�o �o�o+=Oa s2_|_V_���_� ��'�9�K�]�o��� ������ɏ�o���� #�5�G�Y�k�}����� ��ş������ C�U�g�y��������� ӯ���	��ڏ?�Q� c�u���������Ͽ� ���)�����n� 0��ϧϹ�������� �%�7�I�[�m�,��� �ߵ����������!� 3�E�W�i�{�:�L�^� ���������/�A� S�e�w���������~� ����+=Oa s�������� ����9K]o� �������/ #/4G/Y/k/}/�/�/ �/�/�/�/�/??� @?d?&�?�?�?�? �?�?�?	OO-O?OQO cOuO4/�O�O�O�O�O �O__)_;_M___q_ 0?�_T?�_x?z_�_o o%o7oIo[omoo�o �o�o�o�O�o�o! 3EWi{��� ��_��_���oA� S�e�w���������я ������o=�O�a� s���������͟ߟ� �����B�l�.� ������ɯۯ���� #�5�G�Y�k�*����� ��ſ׿�����1� C�U�g�&�p�J��Ͼ� ������	��-�?�Q� c�u߇ߙ߽߫�|��� ����)�;�M�_�q� �����xϊϜϮ� ���7�I�[�m���� �������������� 3EWi{��� ��������  �b$������ ��//+/=/O/a/  �/�/�/�/�/�/�/ ??'?9?K?]?o?. @R�?v�?�?�?O #O5OGOYOkO}O�O�O �Or/�O�O�O__1_ C_U_g_y_�_�_�_�_ �?�_�?o�?-o?oQo couo�o�o�o�o�o�o �o(o;M_q �������� ��_4��_X�o��� ����Ǐُ����!� 3�E�W�i�(������ ß՟�����/�A� S�e�$���H���l�n� �����+�=�O�a� s���������z�߿� ��'�9�K�]�oρ� �ϥϷ�v��Ϛ���� ҿ5�G�Y�k�}ߏߡ� �����������̿1� C�U�g�y������ ������	������6� `�"߇����������� ��);M_� ������� %7I[�d�>� ��t����/!/ 3/E/W/i/{/�/�/�/ p�/�/�/??/?A? S?e?w?�?�?�?l~ ��O�+O=OOOaO sO�O�O�O�O�O�O�O _�/'_9_K_]_o_�_ �_�_�_�_�_�_�_o �?�?�?VoO}o�o�o �o�o�o�o�o1 CU_y���� ���	��-�?�Q� c�"o4oFo��joϏ� ���)�;�M�_�q� ������f��ݟ�� �%�7�I�[�m���� ����t�֯������!� 3�E�W�i�{������� ÿտ�����/�A� S�e�wωϛϭϿ��� �����Ư(��L�� s߅ߗߩ߻������� ��'�9�K�]�ρ� ������������� #�5�G�Y��z�<ߞ� `�b�������1 CUgy���n� ���	-?Q cu���j���� �/�)/;/M/_/q/ �/�/�/�/�/�/�/? �%?7?I?[?m??�? �?�?�?�?�?�?�/ �*OTO/{O�O�O�O �O�O�O�O__/_A_ S_?w_�_�_�_�_�_ �_�_oo+o=oOoO XO2O|o�ohO�o�o�o '9K]o� ��d_����� #�5�G�Y�k�}����� `oro�o�o���o�1� C�U�g�y��������� ӟ�����-�?�Q� c�u���������ϯ� ��ď֏�J��q� ��������˿ݿ�� �%�7�I��m�ϑ� �ϵ����������!� 3�E�W��(�:���^� ����������/�A� S�e�w���ZϬ��� ������+�=�O�a� s�������h������� ��'9K]o� ������� #5GYk}�� �������/�� @/g/y/�/�/�/�/ �/�/�/	??-???Q? u?�?�?�?�?�?�? �?OO)O;OMO/nO 0/�OT/VO�O�O�O_ _%_7_I_[_m__�_ �_b?�_�_�_�_o!o 3oEoWoio{o�o�o^O �o�O�o�o�_/A Sew����� ���_�+�=�O�a� s���������͏ߏ� �o�o�o�H�
o��� ������ɟ۟���� #�5�G��k�}����� ��ůׯ�����1� C��L�&�p���\��� ӿ���	��-�?�Q� c�uχϙ�X������� ����)�;�M�_�q� �ߕ�T�f�x����߮� �%�7�I�[�m��� �����������!� 3�E�W�i�{������� ��������������>  �ew����� ��+=��a s������� //'/9/K/
. �/R�/�/�/�/�/? #?5?G?Y?k?}?�?N �?�?�?�?�?OO1O COUOgOyO�O�O\/�O �/�O�/	__-_?_Q_ c_u_�_�_�_�_�_�_ �__o)o;oMo_oqo �o�o�o�o�o�o�o�O �O4�O[m� �������!� 3�E�oi�{������� ÏՏ�����/�A�  b�$��HJ���џ �����+�=�O�a� s�����V���ͯ߯� ��'�9�K�]�o��� ��R���v�ؿ꿮�� #�5�G�Y�k�}Ϗϡ� �������Ϩ���1� C�U�g�yߋߝ߯��� ���ߤ��ȿ�<��� c�u��������� ����)�;���_�q� �������������� %7��@��d� P�����! 3EWi{�L�� ����////A/ S/e/w/�/HZl~ �/�??+?=?O?a? s?�?�?�?�?�?�?� OO'O9OKO]OoO�O �O�O�O�O�O�O�/�/ �/2_�/Y_k_}_�_�_ �_�_�_�_�_oo1o �?Uogoyo�o�o�o�o �o�o�o	-?�O _"_�F_���� ���)�;�M�_�q� ��Bo����ˏݏ�� �%�7�I�[�m���� P��t֟����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ 㿢��Ɵ(��O�a� sυϗϩϻ������� ��'�9���]�o߁� �ߥ߷���������� #�5���V��z�<�>� ������������1� C�U�g�y���J߯��� ������	-?Q cu�F�j��� ��);M_q ��������/ /%/7/I/[/m//�/ �/�/�/�/���? 0?�W?i?{?�?�?�? �?�?�?�?OO/O� SOeOwO�O�O�O�O�O �O�O__+_�/4?? X_�_D?�_�_�_�_�_ oo'o9oKo]ooo�o @O�o�o�o�o�o�o #5GYk}<_N_ `_r_��_���1� C�U�g�y��������� ӏ�o��	��-�?�Q� c�u���������ϟ� ���&��M�_�q� ��������˯ݯ�� �%��I�[�m���� ����ǿٿ����!� 3����x�:��ϱ� ����������/�A� S�e�w�6��߭߿��� ������+�=�O�a� s��DϦ�h������ ��'�9�K�]�o��� �������������� #5GYk}�� ���������� CUgy���� ���	//-/��Q/ c/u/�/�/�/�/�/�/ �/??)?�J?n? 02?�?�?�?�?�?O O%O7OIO[OmOO>/ �O�O�O�O�O�O_!_ 3_E_W_i_{_:?�_^? �_�_�O�_oo/oAo Soeowo�o�o�o�o�o �O�o+=Oa s������_�_ �_�$��_K�]�o��� ������ɏۏ���� #��oG�Y�k�}����� ��şן������ (��L�v�8������� ӯ���	��-�?�Q� c�u�4�������Ͽ� ���)�;�M�_�q� 0�B�T�f��ϊ���� �%�7�I�[�m�ߑ� �ߵ��߆������!� 3�E�W�i�{���� ����Ϧϸ����A� S�e�w����������� ������=Oa s������� '����
�l.� �������/ #/5/G/Y/k/*|/�/ �/�/�/�/�/??1? C?U?g?y?8�?\�? ��?�?	OO-O?OQO cOuO�O�O�O�O�O�? �O__)_;_M___q_ �_�_�_�_�_�?�_�? o�?7oIo[omoo�o �o�o�o�o�o�o! �OEWi{��� �������_>�  ob�$o&�������я �����+�=�O�a� s�2������͟ߟ� ��'�9�K�]�o�.� ��R���Ư������ #�5�G�Y�k�}����� ��ſ�������1� C�U�g�yϋϝϯ��� ��ʯ�����گ?�Q� c�u߇ߙ߽߫����� ����ֿ;�M�_�q� ������������ ������@�j�,ߑ� ������������! 3EWi(��� ����/A Se$�6�H�Z��~� ��//+/=/O/a/ s/�/�/�/�/z�/�/ ??'?9?K?]?o?�? �?�?�?�?���O�E�$FMR2_�GRP 1ZE�� ��C4  B�� 	� � VOhLS@Fw@ ~EE���B�~A�:{A�L�FZ�!D�`�D��� BT��@�{�ÖM?�  �O��<S@6����B���5�Zf5��ESQ�MA�  �_0[BHT�@JQ@_�33@�TPXSB�<RDx_�]S@@OQ��_�N�_�_RA<�z��<�ڔ=7��<�
;;�*߲<���M8����9k'V8���8���7�?�	8(���_?o �_<ouo`o�o�o�o�'�,B_CFG [9KThB�o/�i�NO 9J
�F0cq hp�lRM�_CHKTYP  )A� A@C@�0+A�ROM~p_MIN\�p�#���p�oP]X,@SSB�c\E TF���%�s���eTP�_DEF_OW � �$AC$�IR�COM�p5��$G�ENOVRD_D�O�v�!b�THR֥v d�dh�_E�NBT� h�RA�VC2C]�w�p �vE� ��o$��Lq2�C�fZ �ȁ�OU5@c9Lkq8fH9�fE<�p�O���d���ԟ��#C�  D+�1���L�\�@OAC�B�gAI�iI����ɀSMT2Cd�։E@�p'��$HO7STC�b1e9I�p���/R@ MC��$?����&�  27.0M�16�  e-�z��� ������h������:�ѿ˳	anonymous>�l�~π�Ϣϴ��"��Q@�� ��+�-��a�B�T�f� xߊ�Ϳ��������� ��K�,�>�P�b�t�� �����������5�� (�:�L��	������� ������� $6 H������������ ��� c�DV hz�������� �
//_q��� m/��/�/�/�/�/7 ?*?<?N?`?�/�� �?�?�?�?�?3/E/W/ i/k?\O�/�O�O�O�O �O?�O�O_"_4_WO �?N_|_�_�_�_�_O O+O�_?_0osOTofo xo�o�o�O�o�o�o�o o]_>Pbt� ��_�_�_��Go (�:�L�^��o������ ��ʏ�o�1�$�6��H�Z���ߡENT �1f��  P�!鏫�  �� ��֟ş������B� �N�)�w���_����� 䯧��˯,���b� %���I���m�ο���� �ǿ(��L��p�3� iϦϕ��ύ��ϱ�� �����G�l�/ߐ�S� ��w��ߛ��߿���2����V��z�=�QUICC0��c�u���1�����&���2�'���v�!ROUTERw�S�e���!PCJOG�����!192.�168.0.10����CAMPRT,��!1 >�%RT��BT� �!Softwa�re Opera�tor Pane�l�{�NAM�E !��!R�OBO0S_C�FG 1e�� ��Aut�o-starte�d�tFTP� ��ޏ����/ #/5/~�Y/k/}/�/� �/F/�/�/�/??1? �pw��|?�/��? �?�?�?�?�/O0OBO TOfO�?O�O�O�O�O �O�O����qOG_ �?�_�_�_�_�_�O�_ oo(o:o]_�_po�o �o�o�o�o__1_C_ Eo6y_Zl~�� eo�����1� D�V�h�z������o�o ���
�M.�@�R� d�v�9�������П� �����*�<�N�`�r� ��Ǐُ���ޯ!�� �&�8���\�n����� ��ǯI�ÿ����"� 4�w������������ ���������Ͽ0�B� T�f�xߛ�߮����� �����K�]�oρσ� t�Ϙ�������� ��(�:�L�o���������������_ERR g&�����PDUSIZ  �q�^���>~$WRD ?e�R��  guestq�dv�����SCD�_GROUP 3�he i{�I�FT$PAO�MP _�SHEDS $�CCOM��TT�P_AUTH 1�i <!i?Pendan���q�n1!KAREL:*����KC//'/��VISION SCET� �/\/m6!�/ �/�/��/�/�/�/7?�? ?m?D?V>�CT_RL j�8�q�
q�FFF�9E3y?P�FR�S:DEFAUL�T�<FANU�C Web Server�:�2R� L^�<YOkO}O�O�O��O��WR_CON�FIG k��?�?��ID�L_CPU_PC�@q�B�S�%P ;BHUMIN\�~)UGNR_IO���2q�	PNPT_�SIM_DO[V�e[STAL_SC�RN[V ��6oQT�PMODNTOL8�We[>ARTY|X%Q�jVy �ENB�W��
SOLNK 1l -o?oQoco�uo�o�obMAST�EZPijUOSL?AVE m�e�RAMCACHE��o�RO�O_CF1G�ocsUO� ~rCMT_OP@8]R
OsYCL�o+u��0_ASG 1n�G>
 �o�� ����*�<�N�`��r��������k�rNU�M1	
rIP��owRTRY_C�NZ+u�Q_UPD1,a� r8pr�o�n� g�� PR�CA_ACC 2�p�  W&j� FD 9� 4�p 6�ŀq��Rᛖ-)�@ 	�@���� � q�̜}�BUF�001 2q�=� iLu0  �u0ihu00x�D�i�u0��Wxi����������������jf�f�!q�p  qpim�iVu�i!�1�B�UQ�b�r���U��������U�����f�f��f�,u0(s�jSf�uu0/_�Exj�f��f�U�f��f��f��f���f���kf�)u0K�)@hu��@r�h9�hUJ��Y��j��y��U������������Uʆ�ن�ꆴ���u0�[�i~�4�@�i;���2���$�)�-�<)�5�h��<�N� `�r���)�~�)�)� ��)¥�)­�)µ�)� ��)�Š)�͠)�ՠ)��ݠR�"��!�SX�)���)������	��	��N0'= �s�h,�	� 5�	�=�	�E�	�M�	��U�	�]�	�e�tp ��l��t�t� �x|����]`Ќ� �ҕ��ҝ��ҥ��ҭ� �ҵ��ҽ���Ű��Ͱ ��հ��ݰ���)��@)��)������3� �+�2�-�2�5�+�F� +�N�+�V�+�^�+�f� +�n��v��~��}� +�䌣��2❢��2� ����2⽢��2�͢�� 2�ݢ+��+����2� ���z���z��� %�z�-�;�z�=�K�z� M�[�z�]�k�\l�{� \|��򅲋Ѝ��ӊ� ���ӊ򭲻ӊ��� ��Ͳ�ӊ�ݲ��2��`2�'����q2r�G 4�<�5\\�<\PS]R}�H�IS�t� ���� 2023-_09-06\+o�������� �:�2);M�Wwk)�8-1�
T7	@;S���JGh	A:{��0:��//'/^�� i�7�k/}/�/�/�/��,ΑZ�	A��� P�/�/|=<k�Y/F? X?j?|?�?�?�?�?�? �??1?O0OBOTOfO xO�O�O�O�O�?	O�O __,_>_P_b_t_�_ �_�O�O�_�_�_oo (o:oLo^opo�jk� w�S/�o�o�o>1  R K@]o]o��dxP����9: c�9`�'�9�K�9/ K/T�������ɏۏ�,Sd� �r� ���#� �_�_~�k�}������� şן����D�V�C� U�g�y���������ӯ ��.��-�?�Q�c� u������������� ��)�;�M�_�qσ� �σop��o�ox��� ��,�>�E�l� ~ߐ�~��|C	���� ���C�G�Y� k�Y�k��ϳ������� ��鏛��"��� ��C� U�׿鿋��������� ����	-d�v�c u������� <N;M_q� �����&8 %/7/I/[/m//�/�/��/�ϐaI_CFG� 2u�� H�
Cycle T�ime�Bus=y�Idl2��min�+.��Up�&�Re�ad7Dow�+8'?�<1�#Co�unt�	Num� �"����<���1�aPROG�"-v������?�?�O!O3OEOWO29�eS�DT_ISOLC�  ���5�6���$J23_DSP_ENB  �K�,�@INC w��M��@A   ?��=���<#��
�A�I:�o  �A_(_��_P_�G�0�GROUP 1xv�K��< P�C��_X_?��?�_��Q�_o!o3o�_ Woio{o�o�@_b[�IN_AUTO � ���J�@POS�REC�C�b71�hK�ANJI_MAS�K�f�jKAREL?MON y�˰?��yRok}���(�.)r�3z�7�C����u�ouCL_L��`NUM�@
��@K�EYLOGGIN�G�`�����E�0L�ANGUAGE ���q���DEFAULT l���LG�!{�:�72��x�@� � 8,�H  �V��'0�������ycO1�;��
�(UT1:\�� ��.�@�W��d�v����������(�Z���LN_DISP |�O48�_|�_!�OCTOL`����Dz�0�A�Av�GBOOK }���dޔ.��ᑮ�X ٌү�����,�<�0��,�N�*�	��ۉ��QmK��aO�A��_B�UFF 2~�K ���235ݿ�� .���17�'�T�K�]� �ρϓ��Ϸ������� ���#�P�G�Y߆��C~��DCS ��9 �B�AK�����%�� ���$��IO 2���� !Z�Q�]�m������� �������!�5�E�W� i�}����������������8�ER_ITM�Nd�ofx�� �����, >Pbt����8�p�;SEV�`�M]7TYP�NU�6/H/Z/��aRST�(���SCRN_F�L 2�F��0� ���/�/�/??(?:?Fk/TP>��O%"M=NGNAM�Dǥq�n��UPS)�GI� �	��E�1_LO�ADPROG �%g:%	T_AR�CWELDG?�MAXUALRM%�,�a���E
B�1'_PR�4�` ��L�@C,����hO����%��ODoPP 2�.�� �ؖ	%/�O �O�O�O_-__Q_<_ u_X_j_�_�_�_�_�_ o�_)ooMo0oBo�o no�o�o�o�o�o�o %[Fj� �������3� �W�B�{���p����� Տ��ʏ���/��S� e�H���t�������� Ο��+�=� �a�L� ��h�z�����߯ʯ�����9�$�]�HDBGDEF �YE���eOu�_LDXD�ISA�0f;6�ME�MO_AP�0E {?g;
 �� F������/�A�S��e�@FRQ_CF�G �YG��AM F�@���H�<�ԃd%h���yϋ��B��YKL��*�/� **: (�H��-���H�S�e� �߉ߛ��߿�����J� YE'� �N�<�R�`�,(�ߥ������ �����*��N�5�r� ��k�����������~JISC 1�g9� �P�JL���`�K���� _M?STR ����SCD 1�ֽ� �/�S>wb� ������// =/(/M/s/^/�/�/�/ �/�/�/?�/ ?9?$? ]?H?�?l?�?�?�?�? �?�?�?#OOGO2OkO VOhO�O�O�O�O�O�O _�O_C_._g_R_�_ v_�_�_�_�_�_	o�_ -ooQo<ouo`o�o�o �o�o�o�o�o;��MJPT��1���8s{�w^sMI�R 1����p ��L���.s< ��?O��.q?y3�\�N��  ����P���.���©� &��5C��o.q���~ �+yH��@�b���v� ��Ə珺����ҏ D�b�4�^���b����� П��؟�+y����L� ^�����g�q���ͯ k�ů�����K�-� ~�����5�W�ɿ���� ׿ϯ��G�-�?�a� c�q�����g�yϛ�� ����U�;�]ߋ�q� ���ߣϵ���߽� ?���3�=��a��� ����������J�\� �����e�w����i� ��������I+�| ��3U����� �E+=_��o^pKdq�j{ � �\rLTARkM_��ju�p��xtop/$^pME�TPU  .r��]qNDSP?_ADCOL3%��>.CMNTT/ �G%FNp t/E'FS�TLI�/�'MST ���/xs� ?|
4G%POSCF�'=.PRPMs/9[STR 1�j}4�q<#�
�16q�5�? �7�?�?�?�?�?�?�? .OO"OdOFOXO�O|O��O�O�O�O_�AG!S�ING_CHK � �/$MODAQ��jy��@U�DEV 	jz	�MC:t\HSI�ZE3 ��@UTA�SK %jz%$�12345678�9 �_�U>WTRI�fp�j{ lju% �8oh+oloOm�t�S�YP�Q{uVT?SE�M_INF 1���XQ`)AT&FV0E0uo��m)�aE0V1�&A3&B1&D�2&S0&C1S�0=�m)ATZ�o@'tHDl�a`o�#xA������ �oC��o ,��P������� �֏?�Q�8�u�(�:� ��^�p��������)� `�M�����>����� ˯ݯ�����Ɵ؟� [���������h�ٿ �������3����i� �.�@�����v���� ���пA���e�L߉� ��NϿ�rτϖϨ�� ��=�O��s�&ߗ�R��������m_NIT�OR� G ?�[ �  	EXESC1�"3�2:�3:�E4:�5:�`<�7:�8:�9:�5�ҟ� 9��E��Q��]�� i��u������T���2��2��2��U2��2��2��2��U2��223���3��3E�@QR_G�RP_SV 1���k (�A?�=��!4 �{ ����Q_D��^�IO/N_DBJP�N]�!_  �hPcX�? �� �L��20� eV��N   k=ƀ�L�cY-ud1�U�����aPL_NAM�E !e���!Defaul�t Person�ality (from FD)�RR2� 1��L�XL�x<�hP d�"J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j?@|?�?�?�?�?aS2F/ �?OO%O7OIO[OmOO�OaR<�?�O�O�O �O__'_9_K_]_o_��_��F�O�^
�_�_�P�_oo/o AoSoeowo�o�o�o�o �o�o�o�_�_O as������ ���'�9�K�]�, >������ɏۏ��� �#�5�G�Y�k�}�������� H�6� H�b H\�<��   �����dܓĐ�#��E� S�Ő���=����������� ��ٯϯ ����5�W�� hz������	`ï�Ͽῠ�:�o�A!"��%�7� �A�  Lɨ�'Ttw.����k��e~� �G��hȟ���� ���������
�C���R� 1��u���@ � ������ @D� M ��?��Ӂ�?�����A��6Ez�  �ј��;�	�l��	 ��@� c0vw�� ����� � � ���� J��K� ��J˷�J�� �J�4�JR�<(�7'��d��� @�S�@�;�fA6A���A1UA���X@�O��=�N���f������T;f��X����E��*]��  �5��>�]���ҘM�� �?����#�������6�w�(� ��>�=���P�H�Ҭu�u�(y���u��Ï�5߫�N�	�'� � ���I� �  y�Y�L�:�È��?È=���Q��� <���� � �� _H��?����I�p�~��e��z��@!��p@�a�@��@ھ�@��C��CR� �� ��B��C��d�@�7�����~3����K�L�����I�@�m�D�՚��������(
%Y:�a�  =�x?��ffd�K/]/� ���/�+R�8Y �/�*>��=��I�� �&��6)������_�>���A!E�<2��!<"7�<L���<`N<D?��<��,-�j?�y/�����"I�?offf?m?&�0�q�@T싹1?��`?Uȩ?X��1W	�1���� ���?��O�7��|/QO <OuO`O�O�O�O�O�O`�O�O_W�5F�  _S__w_�?�_Ij_��_fXHmN H[��YG� F���_oo
oCo.ogo Ro�ovo�o�o�o�o�e t}�o`��_T�_{ �o����t?����/��S�>�w�b� U��Uɲ�Cq�֏m���������D�,/�W	ç��®���+BH� �� T���� ������@I��Y�@n�@���@: @l���?٧]�� ���%�n��߱���=��=D��������@�oA��&{C/� @��U���+J8���
H��>��=3H��_E�� F�6�G���E�A5F�?ĮE��m�����fG��E���+E��E�X����>\��G�ZE�M�F�lD�
�� ����
���.��R�=� v�a�������п���� ߿��<�'�L�r�]� �ρϺϥ�������� ��8�#�\�G߀�kߤ� �ߴ���������"�� F�1�j�U�g����� ����������B�-� f�Q���u��������� ����,P;t _��������:%7p+�(�-�4�t-1�y��]3�ϩ�<���4 �{�����0+#����jb/+/1E�䴛|�0G+E)�/@s/�/�/�/�,.uPe2	P�.q(?{4? ^?I?�?m9F ��?�?@�?�?�?�?�?��$O OLO7OpO[O�O;?�O�O�O�Le�O�O1_`_A_g_U_1)m_�_�_�_�_�_�_j  2 H�6���H�@",c\���B�������Bȓ���A��@��so��w��o�o�o�o�o1v#o5oP,>P`|���T%�����Aotc��
 `��� ���&�8�J�\�n�`������#�rr����H-��$MR�_CABLE 2}��( V`�2T0aa@3 ?0w��ab��{�?`�B?`C �3!OM��`B���3"�z��3!E�33&����J`�N`B��S`�O
�v7��^E!��3 G��@*���X�j�Z`��J`CW`9-��u�7�돒c���gm�Y�����*!���S` �C�/�7� 7��E!�2vouD�r������ Z�+u�M�_�į��ͯ �����ݯ�T�O�%� q�I�[����ɿ7��!���(�:�1(�iϸ{ύ�1(*��*�* ݃OM �����HV3"��]%% 2345678901�ς�� ����3  � 4ba�3!
כ��not sen�t ��?�W�%�TESTFEC_SALGRPg0*"bad�ԈqF�
��0�0k~h������1(9UD1:�\mainten�ances.xm�l�_�  �z��DEFAUL�T�l݂GRP 2=���  p�tg�3%  �%1s�t mechan�ical che�ck�3!�������U� �j7��I�[�m��3"��co�ntroller ��������T(���`!3E��M��,m3""8�3 ���U������P
C��3�W����������C��ge��. b?attery�G/�U	tI/[/m//��/��Supply greasQ,�/����#<��!�/�U8/??1?C?�U?���cabl�/�/�?,(
�/�?�? �?OO�����?�?��?�O�O�O�O�O�%@$�O_Ը׿4_  �OY_k_}_�_�_�O�_ _&_8_�_o1oCoUo go�_�o�_�_�_�o�o �o	jo�oQ�o@ �o�����0� �f;��_�q����� ���ˏ�,��P�%� 7�I�[�m�������� ǟ�����!�3��� W�������ܟ��ïկ ���H��l�~�S��� w�����������2� D��h�=�O�a�sυ� Կ����
������ '�9�Kߚ�o߾����� ����������N߶�5� ��$��}������ �����J��n�C�U� g�y����������� 4�	-?Q��u ���������� f;��q�� ����,/Pb 7/�[/m//�/�/� �//(/�/L/!?3?E? W?i?�/�?�/�/ ?�? �?�?OO/O~?SO�? �?�?�O�O�O�O�O2O �O_hO_�Oa_s_�_ �_�_�O�_�_._oR_ 'o9oKo]ooo�_�o�_ �_�oo�o�o#5�l�b	 TCp� ��o������ !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w����������џ�����+�=� � ��a?�  @�a �x�������fd�ɯۯ�h;*�** �a�f ��?�A�S�e�'������������o�c$� ¿�"�4���X�j�|� ƿؿ�P�������D� �0�B�Tߞϰ�ߜ� ����
ߔ�����d� v߈�&�t���Z�������*�<�j�$M�R_HIST 2���e;�� 
 �\�b$ 2345?678901K�S���J�9�o���� s����o(���� ^p�9K��� � �$6�Z ~�G�k��� /�2/D/�h//�/�/U/�/ �SKCF�MAP  �e�>���z �z �/�%ONREL  z$;��!� ��"EXCFENB�%7
�#�%>1FNC�E?74JOGOVL�IM%7d;�0�"K�EY%7�5�5_�PAN$8�2�2�"R�UN�<�;SFSPDTYPe805�#�SIGN%?74T1�MOT�?41�"_�CE_GRP 1��e�#C�[p�� �Oz#|O�O&D�O�O�O __�O>_�ON_t_+_ �_O_�_�_�_�_o�_ (o�_Lo^oEo�o9o�o �o�o�o�o�o�o6��k�!QZ_EDI�T"D�'CTCOM_CFG 1��-aH5��� 
vq__ARC_B2%E�p9T_MN_MO�DE"F�P9UA�P_CPL�T4N�OCHECK ?��+ �/  S�e�w���������я �����+�=�O�a��;NO_WAITc_L!GkwV@NT~q���+�ez#��_7ERR`A2��)�!���
��.���1S��e����pOᓫ�|� FX+��z!<�0�� ?���Я���0��ڒPARAM:⒬�+�O����S�>��!p��� =  ����������ۿ�ɿ ��#�5��Y�k�G�=���ϯ�B���BODRDSP�s$FP8�OFFSET_C�ARap$�	�DIS���S_A�pAR�K"GlyOPEN_FILE5�$A�qlv��pOPTION_�IO�?�1��M_P�RG %�*%$�*����i�WOU�-�fGP���	��z$��   0 � z$#���#�	 чx(#�z&������RG_DSBL'  3��!̚�����RIENTTO�$0z!C�0�!A�)���UT_SIM�_D���"P���V~��LCT ����hr�q�z%d��_�PEX �8�+�RA-T � dP5+�ПUP ���|�"�������z �􀕕z z 2�1����$�2_C�L��XL�x��%���+=Oa s������� '9K]o�z'2����� 
//./@/R/ã�|/ �/�/�/�/�/�/�/? ?0?B?�il&k/|>��|?�?ϒP�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�?�? _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo �O�OTofoxo�o�o�o �o�o�o�o,>`Pb��Co=����}!�����~�� ��}�}��W�B�{�.�9�p���������ҏ ؏���n���<�K�I�p�	`��~�������:�o����ҟ�|����A�  ��i�'��.�����a��e?b �������e��� q��������˯��������Os�1� ��� � ��>l�@ �]��~G� @D�  Z�?�`�F�?��b���?D�  Ez|�Y5~�  ;�	lr��	 �@�� 0�g�h��� �V�� � � �в���H0#H���G�9G����G�	{Gkf����S��,���C���\���D	�? D@ D��	�������  �O5��>t�[�ù�b�tφ� B��Bp{�!����O�^�#�8��ρ а�������Y�6���:�(:��:��]�T���p��	'� � ���I� �  ����=��������^��� �<��� �� � � *�^��u�^��5���N��\�&���t�?����C��C����B�[���J���i0Z���@�����������A�������
�@�� 2�v���_�\�G���k����������������:�!���x?��ff%�"�� [�Wi��8���
>���n���I� �X����������$��>���
�<2��!<"7�<L���<`N<D?��<��,�/�>`���
�?offf?2�?&lޗ�@T�~?��`?Uȩ?Xǎ�9��gs��� b��`��P��A/ /:/%/^/I/�/m/�/ �/�/�/�/�/?�/6?����/?�?+8Hm�N H[���G�� F���?�?�? �?O�?,OOPO;OtO _OqO�O�E9��M�O%� S?_w?@_�Od_v_�_ �_9�_�_[_�_�_oo<o'o���fb��wkC6o�o2o�o�m?���o�o	�o��Kçs��sm��H��E���Z�d��`��a�q@I܊�@�n�@��@�: @l��?�٧]j ���%�n�������=�=D��ɺ�p��@��oA�&{C/� @�U�� �+J8���
H��>��=�3H��_
� �F�6�G���E�A5F�ğ�E��2�D����fG��E���+E��E�X�Z�D�>\�G��ZE�M�F?�lD�
[��� iϏ���ޏ��;� &�_�J�\��������� ݟȟ���7�"�[� F��j�����ǯ��į ���!��E�0�i�T� y�����ÿ���ҿ� ��/��,�e�Pω�t� �Ϙ��ϼ������+� �O�:�s�^ߗ߂ߔ� �߸������ �9�$� I�o�Z��~�����@��������5��r(�q�4�9����<j�"�3�ϩZ�l��q4 �{�����q��0+#�������jb����1E����|[
	J8�n\���EP*P��A�O�@��#G2 �MT� x����r$�� /�5/ /Y/ �O�/z/�/�,e�/�/�/�/0?,??�A)2?D?�z?h?�?�?�?�:  �2 H�6�vHY��3\��vBoaLcao`B�XpWpA�p@so8OJO\OnO�O�O�M�CP/�O�O�O_T_%\�vN$�p��p�A4T�3�u
 %__�_�_�_�_ �_�_�_o!o3oEoWo�io�z7R����H�-��$PARA�M_MENU ?�
� � MNU�TOOLNUM[-1�w�`F�`�`��iAWEPC�R�`.$INCH�_RATE�`S�HELL_CFG�.$JOB_BA�Sp WVW�PR.$CENTER_RIr�`$t�AZIMUTH �OPTB�a$tE�LEVATION� TC�a$tDW�qTYPE SN�qARCLINK�_AT(pSTAT�US�c�y__VA�LUq�`LEP>�a.$WP_�`�b ��|�����$��6�_�Z�l�~����aS�SREL_ID � ����US�E_PROG �%�j%�����CC�RTƄ��c�_H�OST !�j! �]��T� '�y��@�R�{����_T�IMEOU$��g � �`GDEBU�Gƀ�k��GINP?_FLMSKޟ��TR��PG�p e ���OL�CH�(�yr�k�@���� ү������C�>�P� b���������ӿο� ���(�:�c�^�p� �ϫϦϸ������� ߀�;�6�H�Z߃��W�ORD ?	�k
? 	RS;�Z�PN�q[MA�Ip��SUNq��T�E��ZSTYL5r��COLX�
�Z�L�  �U��0�d�TRACECTL 1�
��a � �� ��M�DT �Q�
��d�D� � � �5P��@��!��"��TQ��p���MP��TIP������	��
����� �ࡐ��7P�㐾䐪��������R����� � � � � �Ȁ�U � � � �U � � � �� � ����R�����㖾���U���������U�N��V��^��f�U�n��v��~����U������������U��������������������lQ������������� ����'�9�K�]�o� ���������������� #5GYk}� ������ 1����//)/ ;/M/_/q/�/�/�/�/��/�/�/?I�LEpȁ]P�`�=�I�?_UP ��[PqY��q ���NQY��}d�bG_zj?�zj�0�&�_DEFSPD ��k{2Ђ  Т`�INPTRL ɵ���a8dU�QPE�_CONFIP�X��̈́}a_0$�LIDS���g0	g�LLB 1�X��P�dTB�  B4Vc}fn�Obljio��eW_ << ρ?��k�o�o�o �o �o6Nl Rd�����ZZo��=�4�a��fQ��C�����ď
eGRP� 1�;l�,�@��  �[�0 � A?x�D P��DV�C2���k��E�d-�=��Q_0����o&aY�#´��r�[�B�����������П����_a>'oY>a����K�]�G� =N�=R�b���^��� ѯ�����z��=� �xM�s�^�  Dz����_`
��ɿx�ٿ�� �#��G�2�k�VϏ� zό��ϰ������j��)Q
V7.1�0beta1_d�60B(�A�?\)A�G���F��>��^����F�A���n�f�fF�A�p��AaG��q�q@�����V�0�ߵ��������p@�
�U`� #�5�G�BҢQ���� �z��v�����F�0B�ga���Ru0��e@:�4+�a��QG�@��0�� B{PB���z�BH�����1�0��g��;Q)���x��xR�N�0n��0��R {�w���W�q�dKNOW_M ��1�c+VdSV �����U ��I[m��|�P�_b5�
cMރ��`�V�	BU����3/�CTߞ��?��@ {Q{�{Pr%n/�,�pa+MRރ��T�כּ�
��/�+̍OADB�ANFWD�+cS�Tށ1 1�Y84�Uk�V�l?_V T?f?x?�?�?�?�?�? �?�?;OO,OqOPObO �O�O�O�O�O�O_�O__572@<	!S?_`G�<}_Q_߀3g_y_�_�_574�_�_�_�_575oo1oCo57A6`oro�o�o577�o�o�o�o578*�<57MA 06��ds�WOVLD  �\{,/ȏ72PARNUM  C;���63SCH�y �u
B��P�.3b�UPD��um����U_CMP_��p���/',5ĄER_wCHK҅��,10"�Ϗ�RS� #?N�_MO ?C�_0�~�U_RES_G?0�\{
��]����� ֟���+��0�a�T� ��x���������fP����Я���P��� ��`,�K�P���_`k� �������`��ɿο�� p��υ�Xp(�G�<Lυ�V 1�F�P�	!@[l�F�T?HR_INR� �q��,5d��MASS6�� Z��MN�����MON_QUEUE �\u,6S��U�TNɀU�N
�3�J�ENDO�m�i��EXEx�iՎ�BE�w�Y�J�OPTIO�V�v�M�PROGR�AM %-�%�LІ�1�K�TASK�_I�t��OCFG� �-��!�T�D�ATA��]�~��2%�������� ���/�A�S�e�w�"������������INFO�ǡ�<ԍ�* <N`r���� ���&8J@\n������ȡ�c ��S�I�K_W���]��ENB��p�[Q&2/(G�W�2�� X,�		�=���&j/�%�!$N0���)�)���_EDIT �]��/�/P�WERFL�خ�23�RGADJ �^�*A�  55?���A5��6M���\u��?�  Bz3W��<�!����%n�?8�/W3�2Y�c7�	HD�l�ǩ��p1?� Ax�ɻt$F*%@/'B **:0B��#O�5CQM\ujBeE��AoI���?�O]M �MmOO�O�O�O/_�O �O__!_�_E_W_�_ {_�_o�_�_�_�_�_ soo/o]oSoeo�o�o �o�o�o�oK�o5 +=�as��� #��������9� K�y�o���������� ۏ�g��#�Q�G�Y� ӟ}�������ş?�� ��)��1���U�g��� �������ӯ���	� ��-�?�m�c�u�￙� ��ٿϿῦ�	p�z� �0hϡό�I��C����ϋ��&�S7PREOF �c:�0�0�
5IORITY����&�1MPDSaP��:���UT?�|C6ODUCT<���*)��6OG�_TG0A��*���HIBIT_DO�	8�TOENT �1��+ (!?AF_INE��^�~�7!tcpi�>��!ud���?!icm��>���XY\3��,��1)� =A�/��0��X�;�G���k� ������������&@8\C��*��\3�c9��?���3�>lK�7�=G/�GL�9�4��8�>A~�2,  �YЀ�����5�6)Z)�
//./�3��ENHANCOE ճ�2A�Ad(�/u%��B��J��\�11PORT�_NUM���0�x�1_CART�REP���S2SK�STA��+�SLGmS[�����3��0Unothing�/s?�?�?�<Y?��?�?�?��61TEM�P ����?8���0_a_seiban��bO��rO�O�O �O�O�O�O_�O(__ %_^_I_�_m_�_�_�_ �_�_ o�_$ooHo3o loWo�o{o�o�o�o�o �o�o2BhS �w������ �.��R�=�v�a��� ����Џ���ߏ���<�'�`�O61VER�SI������ �disable��"KSAVE ����	2670/H755J�]����!~/�����/� 	�S���:�I�|��e@��¯ԯ���J����.�9����_�� 1���|�T��������;�URGEbM B �$���WFİ ��h"��WW�崖���*WRUP_DE?LAY �>ص�R_HOT %�_Ƹ�}/e���R_NORMALD���T�<��x�SEMI�Ϯ�|��9�QSKIPd�	ܺ'u�x[�2�W�V� h�z�=�Gš߯י��� ���߹���'�M�_� q�7��������� ����7�I�[�!�� m��������������� !3EU{i����G��$RBT�IF�
<RCVT�MOU75��� DCRd���� �I�B����C4�BJ���@�.�@�I��*2T�=��]�S]¶f�� �h�����`?�B@�=ߍ��� <2�!<�"7�<L��<�`N<D��<��,�V���- /)/;/M/_/ q/�/�/�/�/�/�/�/���RDIO_TYPE  k���/�EDPROT_C_FG ��26��BHͳEE9
ѻ2�W; �8� j0�?�:��?��?�? OM�?KO��rO�ߓO ��O�O�O�O�O_�O 5_CWaOf_�-_�_}_ �_�_�_�_�_�_�_1o S_Xow_yoo�o�o�o �o�o�o�o=oBao u����� ���9>�]�� _���������ݏˏ� #�(�:���[����m� ������ٟǟ���$� C��W�E�{�i����� ï��ӯ	�/� ��G7?INT 2�Gɔ1=�AG;� ^�p��2���
Hf�0  ��Ȼ��ٯ����� B�0�f�L�vϜϊ��� ����������>�,� b�t�Zߘ߆߼ߪ��� ������:�(�^�p� V������������� �6��EFPO�S1 1�9  x�)c3�� ������*�w�����$ H��l�+� �a���2D ��+�w�K� o���./�R/� v//�/�/G/Y/�/�/ �/?�/<?�/`?�/]? �?1?�?U?�?y?OO �?�?�?\OGO�OO�O ?O�OcO�O�O�O"_�O F_�Oj_|__)_c_�_ �_�_�_o�_0o�_-o foo�o%o�oIo�o�o o�o�o,P�ot �3��i�� ��:�L���3��� ���S�܏w� ����� 6�яZ���~������ O�a������ ���D� ߟh��e���9�¯]� 毁�
����ɯ�d� O���#���G�пk�Ϳ ϡ�*�ſN��rτ� �1�k��Ϸ��ϋ�߀��8���5�n��Z�2 1�f��"�\��� �����"��F���C� |���;���_���� �����B�-�f���� %���I�������� ,��P����I� ��i��� L�p�/�S ew�/�6/�Z/ �~//{/�/O/�/s/ �/�/ ?�/�/�/?z? e?�?9?�?]?�?�?�? O�?@O�?dO�?�O#O 5OGO�O�O�O_�O*_ �ON_�OK_�__�_C_ �_g_�_�_�_�_�_Jo 5ono	o�o-o�oQo�o �o�o�o4�oX�o Q���q� ����T��x�� ��7���[�m����� �>�ُb�����!��� ��W���{����(�ß ՟�!���m���A�ʯ e���$���H���l����v߈�3 1��=�O�����+� 1�O��s��pϩ�D� ��h��ό�߰����� �o�Zߓ�.߷�R��� v�����5���Y��� }��*�<�v������� �����C���@�y�� ��8���\��������� ��?*c���"� F��|�)� M��F��� f��/�/I/� m//�/,/�/P/b/t/ �/?�/3?�/W?�/{? ?x?�?L?�?p?�?�? O�?�?�?OwObO�O 6O�OZO�O~O�O_�O =_�Oa_�O�_ _2_D_ ~_�_�_o�_'o�_Ko �_Ho�oo�o@o�odo �o�o�o�o�oG2k �*�N��� ��1��U���� N�����ӏn������ ���Q��u����4�x������4 1��� j�|���4��X�^�|� ���;���֯q����� ���B�ݯ��;��� ����[���ϣ�� >�ٿb�����!Ϫ�E� W�iϣ����(���L� ��p��mߦ�A���e� �߉��߿����l� W��+��O���s��� ���2���V���z�� '�9�s��������� ��@��=v�5 �Y�}���< '`���C� �y/�&/�J/� �	/C/�/�/�/c/�/ �/?�/?F?�/j?? �?)?�?M?_?q?�?O �?0O�?TO�?xOOuO �OIO�OmO�O�O_�O �O�O_t___�_3_�_ W_�_{_�_o�_:o�_ ^o�_�oo/oAo{o�o �o �o$�oH�oE ~�=�a�П�5 1�ퟗ� �a�L������D�͏ h�ʏ���'�K�� o�
��.�h�ɟ��� �����5�П2�k�� ��*���N�ׯr����� Я1��U��y���� 8���ӿn�����϶� ?�ڿ���8ϙτϽ� X���|�ߠ��;��� _��σ�ߧ�B�T�f� �����%���I���m� �j��>���b���� �������i�T��� (���L���p����� /��S��w$6 p�����= �:s�2�V �z���9/$/]/ ��//�/@/�/�/v/ �/�/#?�/G?�/�/? @?�?�?�?`?�?�?O �?
OCO�?gOO�O&O �OJO\OnO�O	_�O-_ �OQ_�Ou__r_�_F_��_j_�_�_o��6 1���_�_o�o yo�o�_�oqo�o�o�o 0�oT�ox�7 I[�����>� �b��_���3���W� ��{������Ï��^� I������A�ʟe�ǟ  ���$���H��l�� �+�e�Ư��ꯅ�� ��2�ͯ/�h����'� ��K�Կo�����Ϳ.� �R��v�Ϛ�5ϗ� ��k��Ϗ�߳�<��� ����5ߖ߁ߺ�U��� y�����8���\��� ����?�Q�c���� ��"���F���j��g� ��;���_������� ����fQ�%� I�m��,� P�t!3m� ���/�:/�7/ p//�///�/S/�/w/ �/�/�/6?!?Z?�/~? ?�?=?�?�?s?�?�?� O�?DO*o<d7 1�Go�?O=O�O�O�O �?_�O'_�O$_]_�O �__�_@_�_d_v_�_ �_#ooGo�_koo�o *o�o�o`o�o�o�o 1�o�o�o*�v� J�n���-�� Q��u����4�F�X� ���ޏ���;�֏_� ��\���0���T�ݟx� ���������[�F�� ���>�ǯb�į���� !���E��i���(� b�ÿ��翂�Ϧ�/� ʿ,�e� ω�$ϭ�H� ��l�~ϐ���+��O� ��s�ߗ�2ߔ���h� �ߌ���9������� 2��~��R���v��� ����5���Y���}�� ��<�N�`������� ��C��gd�8 �\��	��� cN�"�F� j�/�)/�M/�xq/WOiD8 1�tO /0/j/�/�/?/0? �/T?�/Q?�?%?�?I? �?m?�?�?�?�?�?PO ;OtOO�O3O�OWO�O �O�O_�O:_�O^_�O __W_�_�_�_w_ o �_$o�_!oZo�_~oo �o=o�oaoso�o�o  D�oh�'� �]��
��.�� ��'���s���G�Џ k�􏏏�*�ŏN�� r����1�C�U���� ۟���8�ӟ\���Y� ��-���Q�گu����� ������X�C�|���� ;�Ŀ_�������Ϲ� B�ݿf���%�_��� �����ߣ�,���)� b��φ�!ߪ�E���i� {ߍ���(��L���p� ��/����e���� ���6�������/��� {���O���s������� 2��V��z��/��$MASK 1ꊡ+����XNO  ���?MOTE  �$�G_CFG ��N��PL_RGANGJ?�%��OWER �%���SM_DRYPRG %�)��%K��TAR�T �	*UME_PRO��e/��$_EXEC_E_NB  ?��GSPD> � �(��(TDB�/�*R�M�/�(IA_OP�TION����!_AIRPUR� F*B?.�MT_� T�L2�`1g�o=�";C�?  N?�?��?�?�??1OBOT_ISOLC��>0~zENA_ME F*T/��	OB_CATEG� �O�D�uCORD_NUM� ?�;1�H755  �?�O�OY� PC_TIMEOUT�{ x� S232g�1��# L�TEACH PENDAN!Pc��pT�=JH M�aintenance Cons?�m_?"�_DNo Use�=�__��_�_oo%o�9RN�PO #R�5�6QCH_LA �̋?� 	�aso!OUD1:�ouoR� �VAIL�A5�|�1SR  /;�1��eR_I�NTVAL6��Yp> yV_DA�TA_GRP 2��� D>pP�����y �!��A�/�e�S��� w��������я��� +��O�=�_���s��� ��͟���ߟ��� K�9�o�]��������� ǯ�ۯ���5�#�Y� G�i�k�}�����׿ſ �����/�U�C�y� gϝϋ��ϯ������� �	�?�-�c�Q߇�u���߽߫����$S�AF_DO_PU�LSK�A? ��CS'CANR6�<@�SC�� �`�X�!? �1
�2��A(�Q�U[�? ��� ���������|��#�`5�G�Y�k�HrcE�2��[��d����>	X�Hi @������?��. ��p�_ @3T01n��~�YT D��� ����"4F Xj|�������BoLe��V,/>/F$
*  =iU;�o�Tg!�EqpduE
�t��Di�@�k�Z?  � �+Jk� ��AS��/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_.a����_ �_�_oo)o;oMo_o �_���o�o�o�o�o�o��o	-2qoo0 �"�#�%�-~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N��_r��� ������̯ޯ��� o8�J�\�n������� ��ȿ3auk��� ,�>�P�b�tφϘϪ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{��������(������/�A�S� e�w�������������@��+=��
��T������"�z�	1234�5678�"h!?B!������
���f�� '9K]o��	� �����//(/ :/L/^/p/�/�/�/�/ �/�-��/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO�/�/TOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_3O �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�_�o $6 HZl~���� ���� ��oD�V� h�z�������ԏ� ��
��.�@�R�d�v� 5�������П���� �*�<�N�`�r����� ����̯�����&� 8�J�\�n����������ȿڿ����"����D�V��{ύϟ���
Cz  Bp���   ���2��� }� 6��
���  	���2<�#�5�HG�Y�i���j��� ����������	��-� ?�Q�c�u����� ���������)�;�M� _�q������������� ��%7I[m��� j�k���<� ��  �������
�
�t  ���
"��`�$S�CR_GRP 1��*P3�0 �� ���� ��	 _m�u �k����ǒ�8��������C� ��݌*'����LR M�ate 200i�D 567890��LRMc# 	?LR2D j ��?
1234i%��x�m�� �&_ u��d�d�ӻ����)	�"?%?�7?I?[?k<��#H�u�$yd�?���?�?�?�#�����?(O�?LO�>K� �h��,W&iso  %>�B���!ƗO�B�D�A���O�  @���E�@���@�O ? �E�BH���_�J�F@ F�`8R@_7Od_O_ �_s_�_�_�_�_�_o ��A�AR1oo.o@oRdB�`o�_�o�o�o �o�o�o�o$H3 lW�~ߥz#��w����������A=@ >ճ����@�@U����k�@�'�,�;ϫ���A�@��v΅�?�5ۀ���"�� ��*��z�!M�Y�k�:�h���
����ß��ҟ����Y/k#DEC�LVL  ������"܂A��*SYSTEM*���V9.10214� s�8/21/2�020 A � �`�o�SERV�ENT_T  � $ $S_NAME !���PORT����R�OTO�� ��_S[PD��J�B��̠TRQ  { 
ɣAXISҡ9קϠ 2 �ɣ�DETAIL_ � l $D�ATETI����E�RR_COD(�I�MP_VEL��� 	:�TOQB�A�NGLESB�DI�S��N���G��%$�LIN(� ȤRECҡ ,�����F�MRA�� �2 d��IDX�����ߠ h��$OVER_LI�MI���vɣOC�CURҡ  �-�COUNTE�R��`�SFZN�_CFGҡ 4� $ENABL�(�ST"���FLA�G��DEBUF�R>[�  �J�ҡ � 
$MIN_OVRD��$I��W�{�s����FACE�|�SA}F��MIXED�̸��d�{�ROB���$NE��PPôH�ELL �	� 5$J��BAS�(�RSR_.�  $NUM_�.B� �1w��U29�39�49�59ڕ69�79�8w�	�R�OO��~�CO��O�NLY�p$US�E_AB���A�CKENBA���I}N۰T_CHK��OP_SEL_9����_PU���M_v%�OU��PNS֠����x�9���M3�T�PFWD_KAR�@���.�RE��$�OPTIONX�$�QUE 鿠D;�Y���$CSTOPIg_AL����EX����ь�(�XT��M1ڹ�2��MA��STmY��SO��NB��;DI��TRIFÄ�.@�INI��Mà���NRQ���END���$KEYSWITCH'�<�����HE=�BEATM�o�PERM_LE�?�G�E<�n�U;�F���<�S��DO_H�OM��O����EFaP����G��STL��C��OM)���O�V_MS�ѻ�ET?_IOCMN�Ӕ�������HK>��
 D -Ǳ�3SU'���MP��.��PO��$FOR=C&�WARN�ѧpv��OM� �@?$FUNC� 7ÙU���AR���2��3�4~b�O�L�Lo��!�UN�LO�%��ED�%��p�SNPXw_AS#� 0$��ADDV�X�$S�IZ(�$VAR~w�MULTIP����� Ao �� $�� ��!	&�� ��'�C;�kOFRIF��۰Sl��~	��[NF�OD?BUS_AD�&�د���CM1�DI�A]$DUMMSY1���3�4���SО� � �X�TE���8n�SGL#!TA��  &8�<#'�x� 5 $ STMT��U#PSEG��U!ByW��%$SHOW]%BANi TPO)F��9�0���ȠVC��Gh� 1 $PC�ܰ� ��$FBkP�(S�P��A���%�VD�� g�� � �A0��0�b�$1� �+7� +7� +7� +75�)96)97)98)99
)9A)9B)9} +7�+7r +7F)8� �859@��8O9	 �8i91v9U1�91�91�91�9U1�91�91�91�9�1�9���G592B92�O92\92i92v92��92�92�92�92��92�92�92�92��93(93593B93�O93\93i93v93��93�93�93�93��93�93�93�93��94(94594B94�O94\94i94v94��94�94�94�94��94�94�94�94��95(95595B95�O95\95i95v95��95�95�95�95��95�95�95�95��96(96596B96�O96\96i96v96��96�96�96�96��96�96�96�96��97(97597B97�O97\97i97v97�c�7�97�97�97��97�97�97�97��4ŲVPk�UТG ٠��.�
 �V��� x �$TORu��  �D�M��RΠ��ߔQ_��R��P��G B��S��C=��'�_qU� 2��YSLu�>�� � � 3ǚ
J�$0��^��"VALU3���A���z��FO�ID_L�ֿ�HI��I]$F�ILE_�����$��J�SAϱ� hҐ�E_BL�CKo�#�>!,�D_CPU<�<�
>�����J�x��R  � PW��ثВ��LAc!S�α������RUN_FLGŵ��ɱ��?� ̵걡�걬�Hิ����5T2A�_L}Io  ��G_O��I�P_gEDI�Ҷ T2��,�4��	��7�]���TBC24 � ��̰� ���,�FT�����TDEC̰A��C���M��������TH�S������R��� . ERVE�������������� �X -$:�LEN`��G���:в�RAk�L�N�W_�i�1:њפ2��MO4��S���I��#�㡩�Ք�:о�DE�աLA3CE���CC�#��_MA� ����׎�TCV�/���T !�0�O�E�2���!s�T���!J��A�%M��"��J�0������F�2���� ����6� JK��VK�!��������J�!����JJ�JJ�AAL��1��1�+�
!/�5��b�N1V�b�!��!�L��_Q!
�Q��BCCF� `ҐGROU��?!���!N��CS��RE�QUIR�EBqUj6љ�$T��2��7������ ��� \w f�APPmR��CL!�
$=��N0CLOr�@	S���U	��
��> �n�M���a���'_MG�� C0�p�0	�BRK�	�NOLD�� RTCMO+��
��J+��P3���������PO���X���6 7 �1!���� ��a��!���PATH�����f؟� ��%�� S�CAj��1�INF9�UC�Д��C0KUM(Y������ 	!á�$*�$*:$ �PAYLOA�J{2L��R_AN��e#L��o)k!_){!��R_F2LSHR	Ԩ!LOp$��'#|�'#ACRL_y� �� �W$�H��!��$H�2FLE�X3��J�� P�ϧ�� �
�|409�  :F� X��Щ7�4[�Z���d�v߈�F1�1E"G��@�߻�������RBE�� ��1�C�U�g�y�� )XFT�����6@XX����1��T�W'QX �0Q��D}H���U�H ����0�4�=�+�O��X�j�|���31��! ��������������A1T;F���EL�@��s��J�� ��JE�� CTR�6ATN�Ƒ	v��HAND_�VB!�31��t"� $�PF2���撣SW��~#� $$M� �	����x��|�@�u�vA@Ơ\ �š��A����
A�A���TU��
D�D�P�G����ST����	��N�DY˰. � �t�} ;П'�1�'�!@^'��}T�0�P�P( 1:CLU^g�2�t$ �p�4� �cA��b��ASYIM�#����#���!�_��(�$ ����x/-/?/Q/c#Jj,|*�����)HD_VIds٨b�V_UNK�ؠ�� c�!J���E���,� �%(�L��-���)�/?���S$4,3w��3HRt�i�%zrͱLF0@�DI� ��O�8�rΰ�c& 0`�I�A�#�<@'��'�?@p20�@ϰ �' � �qMEB�At`B�)�T�PT��`�j���dAE0a�oȊ�~�T����� $DUM�MY1:$PS�_9@RF�0�p$���� FLA��Y�P�S��r�$GLB_T�p���j�N1p��x@:qF�( X ���tST�A��S�BR�M21_V���T$SV_ERb� O��@�X�CL��@�A�@O�ɰGLv�EW��) 4��t�$Y!bZ!bW�����!�sAC�"�����U��* �PN�Ѕ�$GI�Jp}$�� q)�ԼФ�+ L��\��S�}$FS�E�֯NEAR�@N@CF<-�@TANC@B"`��JOG�0 �,�0$JOIN�T�Q�P���MSE]T��-  ��E��A�`S�bjp���`��_.� BpU�A�?���LOCK_�FO� �q�BGL�V=sGL��TES�T_XM3 ��EM�Pi��������c$U�0���P2*�����!�+��p��!�)�B�CE����B� $�KAR�AM�TP�DRA��_�V�VE�C�0p�Z�IU!�,�&�HE��TOOL�C��VDREw�I�S3�5��6C6@ASCH|���-��O��rô�30a��SI�#  @$RAIL_BOXE�Q�e�ROBO��?��e�HOWWAR�1����ROLM ��7�a��H�a��*@nvO_F�`!eПHTML5��Оr����w/b�	�Rz�O�20��0k��o 	 ��OUN~�1 d���))��r�a��$PIP��N�P������H@!��� �0CORDED0���� *�XT� ���)ɰ�`O)� 2o D ��OBE� s��P?����?S��qSYS?ADR�qɰj�TCH�p o3 ,�PENҲ*O1A��_����a��ePVWVAE�4 � e����PREV_RTR��$EDIT�V/SHWR�a,� ��B��٠DT��1�'$ a$HEAD�d���A t��KE|�Ѩ�CPSPDX&�JMP\Lᵓ0R��@�5GD1�Ij��SrC^pNE��<qTwTICKC��MM1~'HN"��6 @I�!�e`!_�GP�&��P0STY���LOѝs�"�"��07 t 
�G��%$���=,�S`!$��PY�������P��&SQU�Y��5��ءTERC�n�!a��S�d8 ��8��g�P�g%Q��b�`Oo�b�D@IZ��4������PR%���B�!� PU�aE_�DO2�XSz�KN�AXI<@[&�UR�`�Cr � jd�q�`_��|ET}BQP��Xҕ;0Fҗ�<0A߁Ց��9���)����SRqt9l�0�y�R�z�E �v
Y�r�E�w�C��C �>U3�>UC�>US�PU@j]��PU�\��nYC�_|]C�]L�^�p������SSC�� : �he�DS� `��S�P�jeATA��r�A� �"��ADDR�ES��B�SHIyF�c�_2CHp�fIмa�TU��I�q ;�COUSTO�D�V��I�<���~aC��
��
7V�-AG�'= \*���;0|�1�0IrC��2�Bz��^�Iq�TXSCWREEA>ٰW1TINA{��Мt����~A~b��? T �![�B|Z�7��vJAp{JB�t�RRO��G�{R �q8��UE��$@ ��@���S�|�|RSM� @GU`.�0�S�ͰS_�Ӏs��c�v����~ACx��O��t 2?ǰUE��A�kҶ�@WGMT_�L9�YAzG�Ol�BBL_��9W��G�B �;0�5O���LE�b*�x �b)�RIGH3��BRDmԤaCKG�R��[�T/Z�W�WIDTH�� 7¾�|�����UIj EY~`F�C�z 6 �2��	ABACK�1BΕq�M�FO��LAB(Q?(�M�I����$UR���Ч�S�H	� OD 8��G�_@!�b1�T�R�����C����� �O�aG�E�� x�T�U?��R��BLUM�aF�`GERV����P1�j��FK��@GE�0�@5I LPѥ�B	E�0/a)�?a��Oa�������5��6��7��8ޢ�2b�@1�]tԳ�����S�0EUSR��G �<*�S�U���c��F�O�`��PRI�Amx��m�аTRIP��m�UNDO�H��`0�BE)AEp̀�{@u0 I,�\��AG H0T[ �a�a'�OSr�<�R �@�Û�ӁJ�ߤ� ��c��$8�U١Ӂ�Kl�~ό�٢�%�OSFF����L(��ÉO��"�Je����Ke�GUvPў�8a)׻�SUB�"t�&�RTe��DM�"F��g �3OR��o�RA�U�@p�T�٢U�_���$N |�@�O�WN��$SRC���^0D�����B�MPFI4a}@ESPA�2�p����.!�����TҬ�
 ӁO M`��WO$P��1n�0COP��$r@��_�м�i��p�WA�C��M�#�L����p�5�a P~�rSHADOW^@����_UNSCAp~�㓔��DGD��WEGACc�w��VC P)�ӁQǔ ��@l3$�ER�p,��1����yC� ,�DRIV�6�A_V� O�� 6 �D|�MY_UBY {�4�B6c�l5��0�pb.!��1���P_��4��L#KBM&��$� DEY�EXX �'�t�MUv X&��h�US]�h@˰_�R�q�2���`��1G>�PPACIN�!i0RG��Xn��n��n��i�REF��ac����n�R �`[�Gt�Pr� ��RS��S��x��d��O�	h�:ARE+�SWf _Ag�$ @O���aA�`'��BEl�U.0H������HK32Tu��?���A$�ppEA�� zL�3�'��MwRCVӁU �ʠUO?0M3�C�s	�8�ð�REF��� �����C� ����!�!�1%�f_ ��|g(�xPSi�����1"2��ЄV ��2�����0������0OU�'��&4� �Q�a2��$0�p_p@��S}ca��!D��`UL�pTf(�COG�H�U 0NT#�P41�O5`�[6��[30L��5����5`��7���VIsA_L�]`W ���HD�`Ɛ$JO�g����$Z_�UPL̰ �ZEPW��5�139���_LIM�$EP1I�4� �1�1�q�a���`�%�>6�X� 0}c�Az@` }cCACH��LO!lD�A �I���|���C@MI�cF�A�ETVP�F�+$H�O3���p@COM	MJ�O�O=��G�'��`d3��͡�$ �VP�<p�6R_SIZ��@T�ZR ;X�1<W��n�M]P`ZFAI�0Gl��@AD�Yi�MR1E�$�REWGPU� ���s�ASYNBU=Fs�VRTD�U�TlEQn�OL�`D_���
eW��PC�`TU� �@QD�UECCU�VEM� �ERb�GVIRC�Qe�S|N��Q_DELA�����簶�AG�YR�XYZ��}�W@��h!�d��o`T�IM�af�b���E_GRABB`�Y+�� %�ЄY.�ڒL�AS���PA_GE�WEZ>���sbc_uT@�#���)����I�tX��fb�BG/�V���p�PKq �fXA�'G%IOpN�)��	�H�@�Q:�[���AS�Pr}FN��LEXPv\��ӳ��z�Q��I �S��E���E���Bm��a����]���+��DY�����*�ORDı��°@��"��^ $0TIT��ɰ������VsSFv���_  ���$�[1 UR�SM��`����ADJ�΀�0ZD�a D��AAL�0�PΠ�
BPERI<@��MoSG_Qc$FQ dU[���eBa�b��뇰0�@���@�W�X�S�h�c��� K��CH)�HOL��] �pXVR�d7r�+�T_OVR2�_�ZABC\�e��6��C�
MAc�z�V�S@ f � �$_���|�CTIVz��AIO���FfY�IT
�mDV	�#
mX@��{Q��MàPS�!�� �S����A� ���ALST`Y��A�00��_S���4�c�DCSCH��g Lg�#�w���@ �GÀ@� EPGN�A�C���A"�_F�UN��@���Z&��h���$L���GqZMPCEF\�i���
���f��LN �.�
 ����`]�j $x�Az��CMCM` ECr�C\����P^�? $J��D+Q!�2�+ǚ07Ś0`Ǩ��0�c�UX�a��UXE&���a&� z�<�z����Ɍ����FTF<1!����Y��k D���7p�4��Y@Dp Wl 8cR�PU��$HEIGHYF�?(0ؖ��p|���$m � �S�$B0A���L�SgHIFvS��RV@!F�����+�C�0� \�-4�D��ְ^s�Ӳ UD���CE��V|���SPHERh� n ,00�F�fX�l�r���FA;1���c���u��S�HOT��_��@S�MIPOWERFL �q�c�k� ��WFD�O`� ��G@� 1� ������� L!��_EI�P���c��j!�AFz0E_�$���!'FT��S��w�3!�x����f���7!R'`MA@����������p��������[!OPC3UA\�
J�!TPz0p���yd��!
PM�&�XY��e�?Ⱥ	�f.�!�RDM�V��g|z�!R90�2	�h�#/!
���@�X�i/o/!ReL�PCp/�)8^/>�/!ROS���,��4�/?!
CEF� MT�@?�k�/S?!	2C{�q?��lB?�?!2WA'SRC��m�?�?;!2USB�?��n�?7O!STM��QO�o&O�O���OКtO�M��I
�KL� ?%�� (%�SVCPRG1��OZU2__P3�@_E_P4h_m_P5��_�_P6�_�_P7��_�_P8ooP90o5kT�]oQ
_ �oQ2_�oQZ_�oQ �_�oQ�_%Q�_M Q�_uQ"o�QJo �/Qso�/Q�o�/Q �o=�/Q�oe�/Q�� /Q;��/Qcݏ/Q� �/Q�-�/Q�U�WQ ��O�BG`�O P��� 'Q����1��U�@� y�d�������ӯ���� ���?�*�Q�u�`� ���������̿�� �;�&�_�Jσ�nϧ� �Ϲ��������%�� I�4�m��jߣߎ��� ���������!�E�0��i��J_DEV ����MC:�t��GRP 2���� �@bx 	�� 
 ,�� q��﬒�����9� � 2�o�V���z������� ����#
G.k }��X���� �1U<y` r�����	/� -/�"/c//�/n/�/ �/�/�/�/??�/;? "?_?q?X?�?|?�?�? �?�?F/O%OOIO0O mOTOfO�O�O�O�O�O �O�O!__E_W_>_{_ b_�_�_O�_�_�_o �_/ooSoeoLo�opo �o�o�o�o�o�o+ =$a�_V�N� ������9�K� 2�o�V�������ɏ�� �ԏ�#�zG�Y�@� }�d�������ן���� ��1��U�<�y��� r�����ӯ�<�	��� -�?�&�c�J������� �����ȿڿ���;� "�_�q�Xϕ�쯊��� �������%��I�0� m��fߣߊ������߀����!���W��d �^�	E��y��`��������	�%�	�<.������G��� G�W�e�O���s����� ����� C���- Q?acu���� ��)M; ]������� /�%//I/�p/� 9/�/5/�/�/�/�/�/ !?c/H?�/?{?i?�? �?�?�?�?�?;? O_? �?SOAOwOeO�O�O�O �OO�O7O�O+__O_ =_s_a_�_�O�_�_�_ �_�_�_'ooKo9ooo �_�o�__o�o�o�o�o �o#G�on�o7 �������� aF���y�g����� ����я'�M��]��� Q�?�u�c��������� �#������'�M�;� q�_���ן������� ݯ��#�I�7�m��� ��ӯ]�ǿ���ٿ� ���Eχ�lϫ�5ϟ� ���ϱ������M�2� D������eߛ߉߿� ����%�
�I���=�+� M�O�a�������� !����9�'�I�K� ]������������� ��5#E����� ��k����� 1sX�!�� ����	/K0/o �c/Q/�/u/�/�/�/ �/#/?G/�/;?)?_? M?�?q?�?�?�/�?? �?OO7O%O[OIOO �?�O�OoO�OkO�O_ �O3_!_W_�O~_�OG_ �_�_�_�_�_o�_/o q_Vo�_o�owo�o�o �o�o�oIo.mo�o aO�s��� 5�E�9�'�]�K� ��o����̏����� ���5�#�Y�G�}��� ���m�ןş���� 1��U���|���E��� ��ӯ������-�o� T������u�����Ͽ ���5��,���߿ Mσ�qϧϕ������ 1ϻ�%��5�7�I�� mߣ�����	ߓ����� !��1�3�E�{�ߢ� ��k����������� -����z���S����� ��������[�@� 	s����� �3W�K9o ]����/ �#//G/5/k/Y/{/ �/��//�/�/�/? ?C?1?g?�/�?�?W? y?S?�?�?�?O	O?O �?fO�?/O�O�O�O�O �O�O�O_YO>_}O_ q___�_�_�_�_�_�_ 1_oU_�_Io7omo[o �oo�o�_o�o-o�o !E3iW��o ��o}�y��� A�/�e�����U��� ���я���=�� d���-���������ߟ ͟��W�<�{��o� ]���������ۯ�� �˯�ǯ5�k�Y��� }�����ڿ������ ��1�g�Uϋ�Ϳ�� �{�����	����� -�cߥϊ���S߽߫� ��������kߑ�b� ��;��������� �C�(�g���[���k� ���������� ?� ��3!WEg�{ ������/ SAc���� y��/�+//O/ �v/�/?/a/;/�/�/ �/?�/'?i/N?�/? �?o?�?�?�?�?�?�? A?&Oe?�?YOGO}OkO �O�O�O�OO�O=O�O 1__U_C_y_g_�_�O _�__�_	o�_-oo Qo?ouo�_�o�_eo�o ao�o�o)M�o t�o=����� ��%�gL���� m�����Ǐ��׏��?� $�c��W�E�{�i��� ��ß������՟�� �S�A�w�e���ݟ¯ ���������O� =�s�����ٯc�Ϳ�� �߿���Kύ�r� ��;ϥϓ��Ϸ����� ��S�y�J߉�#�}�k� �ߏ��߳���+��O� ��C���S�y�g��� �����'���	�?� -�O�u�c��������� ������;)K q�����a��� �7y^p' I#�����/ Q6/u�i/W/y/{/ �/�/�/�/)/?M/�/ A?/?e?S?u?w?�?�? ?�?%?�?OO=O+O aOOOqO�?�?�O�?�O �O�O__9_'_]_�O �_�OM_�_I_�_�_�_ o�_5ow_\o�_%o�o }o�o�o�o�o�oOo 4so�ogU�y� ���'�K�?� -�c�Q���u����ҏ 䏛������;�)�_� M���ŏ���s�ݟ˟ ���7�%�[����� ��K�����ٯǯ�� ��3�u�Z���#���{� ����տÿ�;�a�2� q��e�Sω�wϭϛ� �����7���+߽�;� a�O߅�sߩ������ �����'��7�]�K� ���ߨ���q������� ��#��3�Y������ I������������� a�FX1y� ����9]g��$SERV_M�AIL  g�]�COUTPU}TRh }@GRV 2�;  ` (�-<�GSAVEsa�TOP10 2>� d c/ +/=/O/a/s/�/�/�/ �/�/�/�/??'?9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O0�O_��YP�D�FZN_CFG ;�`$���MQGRP 2�WW� ,B �  A�PgD;�� B�P�  B�4#RB21��HELLPR	����nW ok%RSRoo"o [oFoojo�o�o�o�o �o�o�o!E0i�{�~�  ��]r����r� �h ��r�q�x�r2�h d�|�}8��VHKw 1
�[ � r�|�v���ɏď֏� ���0�Y�T�f�x�࡟�������\OMM� �_��RFT?OV_ENBR���P�OW_REG�_UI0�EIMI_OFWDL������Ue�WAIT-� 1�oR��mQ����wTIMQ���į�VAQ��e�_UNcIT,����LCJ�WTRYQ��G�MON_ALIA�S ?e���he�������úm� ���
��ǿ@�R�d� vψ�3ϬϾ������� ���*�<�N�`�߄� �ߨߺ�e������� &���J�\�n���=� �����������"�4� F�X�j���������� o�����0��T fx��G��� ��,>Pb s����y�/ /(/:/�^/p/�/�/ �/Q/�/�/�/ ??�/ 6?H?Z?l??�?�?�? �?�?�?�?O O2ODO �?hOzO�O�O�O[O�O �O�O
_�O_@_R_d_ v_!_�_�_�_�_�_�_ oo*o<oNo�_ro�o �o�o�oeo�o�o �o8J\n�+� ������"�4� F�X��|�������]� Ï�����ɏB�T� f�x���5�����ҟ� �����,�>�P�b�� ��������g���� �(�ӯL�^�p������>��$SMON_�DEFPROG �&������ &*S?YSTEM*��߷�p��?��R�ECALL ?}��� ( �}5�xcopy fr�:\*.* vi�rt:\tmpb�ack#�=>16�9.254.@�1�20:17084� K�T�f�xφ�}6�a"�4�F�Q��������xyzrat?e 124 �ϸ� ��[�m�ߒ� �:�4964 ;�M��������9�s:o�rderfil.dat(ܥ߷�S�e��w��0�mdb: ��>��K����� ���4�-ߪ���`�r��� Ǣ�3���P����� ߪ�����_q�<�߽�6640��K��� ��tpdisc 0�����[m��tpconn 93E ������S/ e/w/���7/�K/�/ �/ ?�&8��/`? r?�?��(?:?L1Q?�?4�?�?
1 �?�? �?ZOlO~O���GO �O�O�OO!A�O�O�O Z_l_~_�O�O5_G_�_ �_�__!_�_�_Voho zo�_�_1oCo�o�o�o //�/�odv�/ �/6�/Q���? ,O��`�r����?(� :��oޏ���'� �\�n�����@�� ڟ��������G�X� j�|�����2�ŏ֯� ����ïT�f�x���o�h92.168�.137.1:18572�oL�ݿ� �o����ʿ[�m�� ����6�H�������� "ϴ���W�i�{ߎϠ� 2�D��������� ����[�m��$� 6�H��������"��� ���d�v�����6����K����� ��$S�NPX_ASG �2���%�  ���%�M  ?��PARAM �%/ �U	;P��PΡ�&  OF�T_KB_CFG�  �+OP�IN_SIM  %���( RVNORDY_DO  ���:QSTP_DSB��~�SR %	 �� &2 ABWE'LD_������TOP_ON_E�RRG�PTN� % ��A	"RING_�PRM�YVCN?T_GP 2��2 x 	zy/�`g/�/�/�/VDN �RP 1u	�  �!%�/�/?#?5?G? n?k?}?�?�?�?�?�? �?�?O4O1OCOUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�_�_�_oo )o;oMo_o�o�o�o�o �o�o�o�o%L I[m���� ����!�3�E�W� i�{�������؏Տ� ����/�A�S�e�w� ��������џ���� �+�=�d�a�s����� ����ͯ߯��*�'� 9�K�]�o��������� ɿ�����#�5�G� Y�k�}Ϗ϶ϳ����� ������1�C�U�|߀yߋߝ߯������"P�RG_COUNT���"��ENB�4/��M$��1�_U�PD 1�T  
���{��� �����������/� X�S�e�w��������� ������0+=O xs������ 'PK]o �������� (/#/5/G/p/k/}/�/ �/�/�/�/ ?�/?? H?C?U?g?�?�?�?�? �?�?�?�? OO-O?O hOcOuO�O�O�O�O�O �O�O__@_;_M___ �_�_�_�_�_�_�_�_�oo%o��_INF�O 1i�9O�q`	 Ho�o�wo�o�i?�̬@�d�7=��?�q*�o B��;c7���o�g>�CP ?�2 A�6~��b�n >���{ �'���Dd�8C���6���X� �b@p�d���ðXD̿�73���W����3���YSDOEBUG	�j��?`�dR�zpSP_PA�SS	�B?�{L_OG ffs�  ?`xEo � �aq`  U�D1:\�tLn�r_MPC�}i�:�L�i���o>bi��SAV �y�a�q�r�;e �SV�T�EM_TIME �1�wt� 0JO�sK�j��ʇ�MEMBK  i�N���N�`�p��X|O�� @p�;cВ���ǜ��d�����q �k@�/�A�S�e���}��������ůׯ� � ��!�3�E�W�i�{�������e��ӿ��� 	��-�?�Q�c�uχ� �ϫϽ���������)�̅SK%�*��9��i�{ߍ߁�1?`j�,�2����A��p�  ֒"���9f(
���^�p�ԟv�;e� ������@����������߀+�@P�b�t�����?`$�� ��������,> Pbt��������(:.�T�1SVGUNSP]D�u '�u�]�2MODE_LI�M ,�恐rY2�f��}XAS�K_OPTION�p-��q�_DI~�pENB  ����u�BC2_GRP 2LՌs�$/̄��C�9#QBC?CFG +��1����p*`�/�o �/�/�/�/�/ ??D? /?h?S?�?w?�?�?�? �?�?
O�?.OO>OdO OO�OsO�O�O�O�O�O _���L _�OS_e_�O B_�_�_�_�_�_q�o /��Po1ooUoCoyo go�o�o�o�o�o�o�o 	?-cQs� �������� �)�_�E�0Ps����� ��ǏE��ُ��!�� E�W�i�7���{����� ՟ß����/��S� A�w�e�������ѯ�� �����=�+�M�O� a�������q�ӿ�� �'ϥ�K�9�[ρ�o� �Ϸ��ϗ�������� 5�#�E�G�Yߏ�}߳� �����������1�� U�C�y�g����� �������ѿ3�E�c� u�������������� )��M;q_ ������� 7%[Ik� ������// !/W/E/{/1��/�/�/ �/�/e/?�/?A?/? e?w?�?W?�?�?�?�? �?�?OOOOO=OsO aO�O�O�O�O�O�O�O __9_'_]_K_m_o_ �_�_�_�_�/�_o#o 5oGo�_koYo{o�o�o �o�o�o�o�o1 UCegy��� ����	�+�Q�?� u�c���������͏Ϗ ���;��_S�e��� ����%�˟��۟�� %�7�I��m�[���� ����ůǯٯ���3� !�W�E�{�i������� տÿ�����-�/� A�w�eϛ�Q������� ��߅�+��;�a�O����o֣��$TBC�SG_GRP 2�o�� � �� 
 ?�  ������� ��(��$�^�H�����Ү���d@� ���?��	 H�BL������B$  C�����	���f��Cz	�Q�AД��333?&ff?7����A����:a� ���ͷ�|�f��DH����@�q�`��t� ����D"w� ����d/
��r� ���u������:Ic	�V3.00��	�lr2dI	�*�}�ҔS �� ��� � �/+��J2®���fG/$%CFoG !o���Y ��K*�u"�x,�,��/�/�* x��/�/�/?	?B?-? f?Q?�?u?�?�?�?�? �?O�?,OO<ObOMO �OqO�O�O�O�O�O�O �O(__L_7_p_�_�� ���_�_�_[_�_�_�_ oo>o)oboMo�o�o �o�owo�o�o�o :�я�_k�oq� ������%�� 5�[�I��m�����Ǐ ��׏ُ�!��E�3� i�W���{���ß��� ՟����5�G��g� ��w�����ѯ����� �+�=�O��_�a�s� ����Ϳ߿�Ͻ�'� �K�9�[�]�oϥϓ� �Ϸ��������!�G� 5�k�Yߏ�}߳ߡ��� �������1��U�C� y�g���Y������� ���	�+�-�?�u�c� �������������� ;)Kq��O �����7 %GI[��� ����/3/!/W/ E/{/i/�/�/�/�/�/ �/�/??A?S?��k? }?;?9?�?�?�?�?O �?OO+OaOsO�OCO �O�O�O�O�O__'_ 9_�O]_K_�_o_�_�_ �_�_�_�_�_#oo3o 5oGo}oko�o�o�o�o �o�o�oC1g U�y����_? ��!��Q�?�a��� u�����Ϗ����� )��M�;�q�_����� ��˟������%�� I�7�m�[�}�����ǯ ���ٯ����!�3� i�W���{�����տÿ ����/��S�A�w� ��3��ϳ�9�o����� ��=�+�M�s�aߗ� �߻�yߋ������� 9�K�]�o�)���� ����������5�#� Y�G�i���}������� ������UC yg������ �����EW/ u�����/� )/;/M/_//�/q/�/ �/�/�/�/??�/7? %?[?I??m?�?�?�? �?�?�?�?!OOEO3O UO{OiO�O�O�O�O�O �O�O�O_A_/_e_S_ �_w_�_�_i�_�_�_ �_+ooOo=o_oaoso �o�o�o�o�o�o'�K9oY~  �p�s �v��r��$TBJOP_�GRP 2"au��  K?��v	�r�s$�|��ip�@�� 0��u  � � � � ��t� @�p�r	 ߐBL  I�C�� D�w�qe�>��n�j�|�<�B�$?����@��?�33C�S� ��a���ǇI�[�}�����;�2������@��?�〱z;���V�A�g�Ȇ〝 ���6��p>�̧�����;��p�A:�?�ff@&?ff?�ff��ޟa� ��u�󄦁���,�:v,���?L����ʐDH�^�d�v�@�33�����>ʐ������8��a퉡�q=�2�D"� ����������=�9�K�9��ݯ﯐� ������חɿ�����  �����?�Y�C�Q�� �ϋ�E����������L@ߙsC��v2����	V3.0�	�lr2d�t*����t�q�ߤ� �E8� EJ� �E\� En@ �E�pE�� E��� E�� E��� E�h E��H E�0 E�� Eϻ��� �E��� E��x E�X F����D�  D��` E��P �E��$��0��;��G��R��^p �Ek��u����І���(��� E���Н�УX 9��IR]�)�q���(�����v��9��՟���tESTPA�RSr��x�p�sHR���ABLE 1%*�ys��t���Q `�������記w�q��	��
�����.��q����8��t��RDI��q-�?�Q�c�u�����O��	%7I[�S���s ��. @Rdv���� ���//*/</N/ `/r/�}� ��r,��) ����~�������������"NUM [ au�q%���p s�t��_CFG &�;/3=��@�pIMEBF_�TT��*5�s��6V�ERr��!�6�3R� 1'� 8$�ߙr�p7A dp�/  O1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_�_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [����������!�3���A_�|1�6@�5��MI__CHAN�7 �5} ��DBGLVڀ��5�5�ᡀETHERAD ?������G�E��x��血ROUT�0!�
!S�q�D�?SNMASK��3>��255.��w�ୟ��џw���OOL�OFS_DI���k�ӉORQCTRL (Kg��O�T>�s���������ͯ ߯���'�9�K�]� o�������=�ƿ������PE_DETA�Iǈ�PGL_C�ONFIG .��9�1��/ce�ll/$CID$/grp1�d�v��ϚϬ�b�:����� ����1���U�g�y� �ߝ߯�>�������	� �-����c�u��� ���L�������)� ;���_�q��������� H�Z���%7I�.}������ �G1ۿ����6 HZl~����� ���/�2/D/V/ h/z/�/�/-/�/�/�/ �/
??�/@?R?d?v? �?�?)?�?�?�?�?O O*O�?NO`OrO�O�O �O7O�O�O�O__&_ �OJ_\_n_�_�_�_�_ E_�_�_�_o"o4o�_ Xojo|o�o�o�oAo�o��o�o0B=���User V�iew R�}}1�234567890s������tX^�2����Yy2fy �o7�I�[�m������`r3�ߏ��� '�9���Z��4Ώ�� ����ɟ۟�L���5��G�Y�k�}����� �¯�66�����@1�C�U���v��7� ����ӿ���	�h�*��8��c�uχϙϫ�������� l�Camera dzZ�#�5�G�Y�k�}�[Eߧ߹���q�����	��-�?�5�   ���ߏ������� �����1�|�U�g� y������������͉ F���1CU�� y�������� 	�������gy ����h��	/ T-/?/Q/c/u/�/. ��[� /�/�/�/?? /?�S?e?w?�/�?�? �?�?�?�?�/��驊? ?OQOcOuO�O�O@?�O �O�O,O__)_;_M_ __O�����O�_�_�_ �_�_o�O)o;oMo�_ qo�o�o�o�o�or_�� Q�bo);M_q o������ �%�7��o�g9�x� ��������ҏy�� ��+�P�b�t�������9�	��00���� 	��-�?��c�u��� .�����ϯ����� ���۩�^�p����� ����_�ܿ� �K�$� 6�H�Z�l�~�%���r� ������� ��$�˿ H�Z�l߷ϐߢߴ��� ���ߑ�˕����6�H� Z�l�~��7ߴ����� #���� �2�D�V��� �J����������� ���� 2D��hz ����i��+Y  2DVh� ������
// ./��"K�z/�/�/ �/�/�/{�/
??g/�@?R?d?v?�?�?A-  E)�?�?�?�? O#O5OGOYOkO}O�K   �?�?�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q����������L  }
A (  �0( 	 �G�5� k�Y���}�����Ïŏ�׏���1��U���J ��/������ 1?�����*�<�C# ��f�x���џ����ү ����O�,�>�P��� t���������ο�� ��]�:�L�^�pς� ��ۿ�������5�� $�6�H�Z�l߳ϐߢ� ����������� �2� y�V�h�z��ߞ���� ������?�Q�.�@�R� ��v������������ ��_�<N`r �������% &8J\��� ������/"/ 4/{X/j/|/��/�/ �/�/�/�/A/?0?B? �/f?x?�?�?�?�?? ?�?OOa?>OPObO tO�O�O�?�O�O�O'O __(_:_L_^_�O�_ �_�_�O�_�_�_ oo8$ok_K�@ FbSo�eowoFcMg1����+frh:\tp�gl\robot�s\lrm200�id�`_mate=_�b.xml3o�o �o%7I[moV������ ����,�>�P�b� t��������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l���}��� ��Ưد���� �2� D�V�h��y�����¿ Կ���
��.�@�R� d�{�uϚϬϾ����� ����*�<�N�`�w� qߖߨߺ���������&�8�J�\�n�h��Q Mo�`<<w �` ?�n� ��n���������/� �G�e�K�]������ ����������3�aoV�$TPG�L_OUTPUT� 1yQyQ ������ ��0BTf x��������//,/>/P/�����f 2345678901u/�/�/�/�/ �/�#oRr/�/?"?4? F?X?�/\?�?�?�?�?�?n:}�?OO,O>O PO�?�?�O�O�O�O�O �OxO�O_(_:_L_^_ �Ol_�_�_�_�_�_t_ �_o$o6oHoZoloo zo�o�o�o�o�o�o�o  2DVh � �������.� @�R�d�v�������� Џ�􏌏��*�<�N� `�r��������̟ޟ �����8�J�\�n����q}�ᶯȯگ����!�@��E�W���� ( 	  Z/��z�����Կ¿�� ��
��R�@�v�d� �ψϾϬ�������� �<�*�`�N�p�r߄��ߨ���h&������ �*��L�^�8��� b*������q������ ��C�U���Y���%�w� ��������	g���? ��+u�a�� ���);G q����S�� ��%/7/�[/m// Y/�/}/�/�/�/I/�/ !?�/?W?i?C?�?�? �/�?�?�?�?OO�? %OSO�?;O�O�O5O�O �O�O�O_eOwO=_O_ �O[_�___q_�_�_+_ �_o�_�_9oKo%ooo �o�_io�oQo�o�o�o �o#5�ok} �����GY� 1��9�g�A�S����� �ӏ��я�����Q�c���)WGL�1.XML!�����$TPOFF_L�IM ��+�������N_SV���  (���P_MON 2��S+�+�2���STRTCHK �3��������VTCOMPAT՘�_�ĖVWVAR �4����ٔ �6� ��������_DEFPRO�G %$�%	�LABWELD_������_DISP�LAY��$�ʢIN�ST_MSK  �� �INU�SERU��LCK�^�%�QUICKM�EN���SCRE桰��`�tpsc�^��������Ұ_ֹSTS���R�ACE_CFG �5������	
?��HNL� 26٪��A���  ��uχϙϫϽ����������ITEM �27a� �%$�12345678�90H�Z�  =<�R�xߊߒ�  !�ߠ۬�\��ߣ�F� �j�*�<��R����� ���ߺ������v�f� x����(���~��� �����>�P�b����� 2Xj��v�� ��L�*� ���� ��6 �Z�5/�P/�`/ �/�/��/ /2/D/�/ h/?:?L?�/p?�/�/ �/|?�?.?�? Od?O �?�?cO�?~O�?�O�O O�O<ONO_rO2_�O B_h_�O�O�O__&_ �_J_�_o.o�_Ro�_ �_�_To�_�o�o�oFo �ojo|o�o`�o� ��o�0�T� x8�J��`��$��� �ȏ,�؏���t�� ������6�������ğ (��L�^�p������ f�x�ܟ�� ��ۯ6� ��Z��,���B���Ư����S'�8-ϔ�ψ  Ҕ� 89���
 �����B�úUD1:�\O�����R_G�RP 195�?� 	 @렚� �˖��Ϻ��������$�;�I��O�s�^�<�߂�?�  ���� ���������,��<� >�P��t������0�����(�	b�<��N���SCB 2:�� �ߚ������������*��U�TORIAL �;��6�u��V_C�ONFIG <���4��2���OUTPUT =��� ���$6 HZl~���� ����$/6/H/ Z/l/~/�/�/�/�/�/ �/�// ?2?D?V?h? z?�?�?�?�?�?�?�? 	?O.O@OROdOvO�O �O�O�O�O�O�O_O *_<_N_`_r_�_�_�_ �_�_�_�_o_&o8o Jo\ono�o�o�o�o�o �o�o�oo"4FX j|������ ��0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ���� P�b�t���������ο ����(��L�^� pςϔϦϸ�������  ��$�5�H�Z�l�~� �ߢߴ����������  �2�C�V�h�z��� ����������
��.� ?�R�d�v��������� ������*;�N `r������ �&8I\n �������� /"/4/EX/j/|/�/ �/�/�/�/�/�/?? 0?A/T?f?x?�?�?�? �?�?�?�?OO,O>O O?bOtO�O�O�O�O�O��O�O__(_:_����Y_k_UQD_ �_9��_�_�_�_oo &o8oJo\ono�o�oEO �o�o�o�o�o"4 FXj|���o� �����0�B�T� f�x��������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϯ����� ����
��.�@�R�d� v߈ߚ߽߬������� ��*�<�N�`�r�� ������������ &�8�J�\�n�����������$TX_SCREEN 1>mU�UP�}�����	-?Q���V������ ��bt!3EW i{����� �//�A/�e/w/ �/�/�/�/6/H/�/? ?+?=?O?�/s?�/�? �?�?�?�?�?h?O�? 9OKO]OoO�O�O
OO �O�O�O�O_#_�OG_ �Ok_}_�_�_�_�_<_��_�$UALRM_MSG ?����� �_��o-o ^oQo�ouo�o�o�o�o��o �o$H�US�EV  
m�zv�RECFG �@����  ���@�  A�q �  Bȶ�
  I��������%� 7�I�[�m�������q�GRP 2A�{; 0��	 ����PI_BBL_N�OTE B�zT��l�������p��DEF�PRO`%
k �(%MAIN OLD_2ꏶ�%< ��v�����ӟ����⟀�-��Q�<�u��F�KEYDATA �1C��Ӏp �w��֏ٯ�¯��!���,(-�T���(�POINT E�R\�^�WEX�ST������P��߿���END��TO�UCHUP�� � ORE INFO8�;�xϊ�qϮϕ� ���������,�>�%��b�I߆ߘ� ���/frh/gu�i/whitehome.png��`����������point��S�e��w���*���arc_strA�E�������'����weldB�]�o�������4���enK������(��touchup��ew��t�����wrgA� ��/��8\ n����E�� �/"/4/�X/j/|/ �/�/�/A/�/�/�/? ?0?B?�/f?x?�?�? �?�?O?�?�?OO,O >O�?POtO�O�O�O�O �O���O�O_ _2_D_ V_]Oz_�_�_�_�_�_ c_�_
oo.o@oRo�_ do�o�o�o�o�o�oqo *<N`�o� �����m�� &�8�J�\�n������ ��ȏڏ�{��"�4� F�X�j���|�����ğ ֟������0�B�T� f�x��������ү� �����,�>�P�b�t� �������ο���Z������πK�]Ϩ�9φϘϧ�,�~���v�POIN�T ER��n�W?ELD_ST������P�O�
�END�P�Q�TOUCHUP|�}ߨ��߳��� ���&��J�1�n�� g������������K�Dwhitehome�C�U�g�y���>Dpoin����������
9>�c_str��I�[m��(	weld9����2 en�Pb�t��'touchup@���/t/��(wrg8 W/i/{/�/�/���/�/ �/�/??�/A?S?e? w?�?�?�?<?�?�?�? OO+O�?OOaOsO�O �O�O8O�O�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o ��_ko}o�o�o�o�o �_�o�o1C�o gy�����b �	��-�?�Q��u� ��������Ϗ^��� �)�;�M�_���� ����˟ݟl���%� 7�I�[��������� ǯٯ�z��!�3�E� W�i���������ÿտ �v���/�A�S�e� w�ϛϭϿ������� ���+�=�O�a�s�����������߼��ݦ������,��3���W�>�{� ��t���������� ��/�A�(�e�L����� ����������  =$asRo��� ��� �'9K ]o����� ���#/5/G/Y/k/ }//�/�/�/�/�/�/ ?�/1?C?U?g?y?�? ?�?�?�?�?�?	O�? -O?OQOcOuO�O�O(O �O�O�O�O__�O;_ M___q_�_�_$_�_�_ �_�_oo%o�_Io[o moo�o�o2o�o�o�o �o!�oEWi{ �������� �/�6S�e�w����� ����N������+� =�̏a�s��������� J�ߟ���'�9�K� ڟo���������ɯX� ����#�5�G�֯k� }�������ſ׿f��� ��1�C�U��yϋ� �ϯ�����b���	�� -�?�Q�c��χߙ߫� ������p���)�;� M�_��߃������h�����p����p����,�>��`�r�L�,^��V ����������!E W>{b���� ���/S: w�p����� //+/=/O/a/p�/ �/�/�/�/�/�/�/? '?9?K?]?o?�/�?�? �?�?�?�?|?O#O5O GOYOkO}OO�O�O�O �O�O�O�O_1_C_U_ g_y__�_�_�_�_�_ �_	o�_-o?oQocouo �oo�o�o�o�o�o �o);M_q�� $������� 7�I�[�m���� ��� Ǐُ����!��E� W�i�{�������ß՟ �����/���S�e� w�������<�ѯ��� ��+���O�a�s��� ������J�߿��� '�9�ȿ]�oρϓϥ� ��F��������#�5� G���k�}ߏߡ߳��� T�������1�C��� g�y��������b� ��	��-�?�Q���u� ����������^���@);M_6�a��6������������, ��7[mT �x�����/ !//E/,/i/{/b/�/ �/�/�/�/�/�/?? A?S?2�w?�?�?�?�? �?���?OO+O=OOO aO�?�O�O�O�O�O�O nO__'_9_K_]_�O �_�_�_�_�_�_�_|_ o#o5oGoYoko�_�o �o�o�o�o�oxo 1CUgy�� ������-�?� Q�c�u��������Ϗ �����)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� ��h?��ǯٯ���� �3�E�W�i�{����� .�ÿտ����Ϭ� A�S�e�wωϛ�*Ͽ� ��������+ߺ�O� a�s߅ߗߩ�8����� ����'��K�]�o� �����F������� �#�5���Y�k�}��� ����B������� 1C��gy��� �P��	-? �cu�����ڦ���������/-�@/R/,&,>?�/6?�/�/ �/�/�/?�/%?7?? [?B??�?x?�?�?�? �?�?O�?3OOWOiO PO�OtO�O�O���O�O __/_A_Pe_w_�_ �_�_�_�_`_�_oo +o=oOo�_so�o�o�o �o�o\o�o'9 K]�o����� �j��#�5�G�Y� �}�������ŏ׏� x���1�C�U�g��� ��������ӟ�t�	� �-�?�Q�c�u���� ����ϯ�󯂯�)� ;�M�_�q� ������� ˿ݿ���O%�7�I� [�m�φ��ϵ����� ����ߞ�3�E�W�i� {ߍ�߱��������� ��/�A�S�e�w�� ��*���������� ��=�O�a�s�����&� ��������'�� K]o���4� ���#�GY k}���B�� �//1/�U/g/y/ �/�/�/>/�/�/�/	?�?-???�A;�>����j?|? �=f?�?�?�6,�O�? �OO�?;OMO4OqOXO �O�O�O�O�O�O_�O %__I_[_B__f_�_ �_�_�_�_�_�_!o3o �Woio{o�o�o�o�/ �o�o�o/A�o ew����N� ���+�=��a�s� ��������͏\��� �'�9�K�ڏo����� ����ɟX�����#� 5�G�Y��}������� ůׯf�����1�C� U��y���������ӿ �t�	��-�?�Q�c� �ϙϫϽ�����p� ��)�;�M�_�q�Ho �ߧ߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{�
������� ��������/AS ew����� ��+=Oas ��&����/ /�9/K/]/o/�/�/ "/�/�/�/�/�/?#? �/G?Y?k?}?�?�?0? �?�?�?�?OO�?CO�UOgOyO�O�O�O����K�������O�O�M�O _2_V,oc_o�_n_�_�_ �_�_�_oo�_;o"o _oqoXo�o|o�o�o�o �o�o�o7I0m T�������� �!�0OE�W�i�{��� ����@�Տ����� /���S�e�w������� <�џ�����+�=� ̟a�s���������J� ߯���'�9�ȯ]� o���������ɿX�� ���#�5�G�ֿk�}� �ϡϳ���T������ �1�C�U���yߋߝ� ������b���	��-� ?�Q���u����� ������)�;�M� _�f������������ ��~�%7I[m ��������z !3EWi{
 �������/ //A/S/e/w//�/�/ �/�/�/�/?�/+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�O�O"O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o�o��!k������Jo\onmFo�o�o|f,��o��o �o-Q8u� n������� )�;�"�_�F���j��� ����ݏď����7� I�[�m�����_��ǟ ٟ����!���E�W� i�{�����.�ïկ� ������A�S�e�w� ������<�ѿ���� �+Ϻ�O�a�sυϗ� ��8���������'� 9���]�o߁ߓߥ߷� F��������#�5��� Y�k�}������T� ������1�C���g� y���������P����� 	-?Q(�u� ������� );M_���� ���l//%/7/ I/[/�/�/�/�/�/ �/�/z/?!?3?E?W? i?�/�?�?�?�?�?�? v?OO/OAOSOeOwO O�O�O�O�O�O�O�O _+_=_O_a_s__�_ �_�_�_�_�_o�_'o 9oKo]ooo�oo�o�o �o�o�o�o�o#5G�Yk}��$UI�_INUSER � ����q��  ���_MENHI�ST 1D�u�  ( ��p��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1�B�T��f�x��)	��63�1/�ŏ׏��� �	'����7��F�X�j��|�r/���edi�t'�LAB_WELD_5�ҟ���|Y.����AB��2�V�h�z�}��-�MA�INE�կ���� �!�+�4įX�j�|���p�����ȿڿ����q������A� S�e�wωϛϞ����� �����ߨ�=�O�a� s߅ߗ�&�8������� ��'��K�]�o�� ���4���������� #�����Y�k�}����� ��B�������1 �.�gy���� ����	-?� cu�����^ �//)/;/M/�q/ �/�/�/�/�/Z/�/? ?%?7?I?[?�/?�? �?�?�?�?h?�?O!O 3OEOWOBT�O�O�O �O�O�O�?__/_A_ S_e_�O�_�_�_�_�_ �_�_�_o+o=oOoao soo�o�o�o�o�o�o �o'9K]o� ������� #�5�G�Y�k�}�hOzO ��ŏ׏�����1� C�U�g�y����,��� ӟ���	����?�Q� c�u�����(���ϯ� �������M�_�q� ������6�˿ݿ�� �%ϴ�I�[�m�ϑ���ώ���$UI_�PANEDATA 1F������  	��}  frh/�cgtp/fle�xdev.stm�?_width=�0&_heigh�t=10	���ic�e=TP&_li�nes=3	�columns=4	��fon�4&_p�age=doub���1�ϑ�)  r3imX߁�  ���� �߼�������Y��(� �L�3�p��i��� ������ ���$�6���Z���� � �z�
  a��������2!�3�E�92d�b�ual��! ��EWi{��F� �����A S:w^�������h�      ��� 6;/M/_/q/�/�/� �/,�/�/??%?7? �/[?m?T?�?x?�?�? �?�?�?O�?3OEO,O iOPO�O�Or��F�� �/�O�O�O_#_5_�O Y_�/}_�_�_�_�_�_ >_�_o�_1ooUogo No�oro�o�o�o�o�o 	�o-?�O�Ou� ����"�f_� )�;�M�_�q������ ��ˏ�����%�� I�[�B��f������� ٟL^�!�3�E�W� i��������ïկ� ������A�(�e�w� ^�������ѿ����ܿ �+��O�6�s���� ������������h� 9߬�]�o߁ߓߥ߷� ����������5�G� .�k�R��v����� �������Ϥ�U�g� y����������F��� 	-?Qc��� n������ );"_F��|�,�>����/!/3/E/W/)�|/��k/ �/�/�/�/�/?i/&? ?J?1?C?�?g?�?�? �?�?�?�?�?"O4OO�XO��B�<��$UI�_POSTYPE�  B�� 	 dO�O�B�QUICKMEN  �K�O�O�@�RESTORE �1GB� � �KO��5_BS0_��m`_�_�_ �_�_�_t_�_oo+o =o�_aoso�o�o�oT_ �o�o�oLo'9K ] ������ ~��#�5�G��oT� f�x����ŏ׏��� ���1�C�U�g�
��� ������ӟ~����� v�(�Q�c�u�����<� ��ϯ�����)�;� M�_�q��~������ ݿ���%�ȿI�[� m�ϑϣ�F�������x����GSCRE�@�?�Mu1�sc*Pu2J�3�J�4J�5J�6J�7rJ�8J�'�TAT�M�� �CB��JUScER,�1�C�ksLӪ��3��4��5��6���7��8�ъ@ND�O_CFG H��K���@PD������Non�e�B��_INFOW 1IB�q��@0%ߌ���z��� �������'�
�K�.� o���d����������L�^�OFFSET L�Iu�����#P ��,>Pb��� ����( UL^������O��/
/:/���UFRAME  ���.�[�RTO?L_ABRT^/Y��v"ENB/p(GR�P 1MY�ACz  A��#�!3� �/�/�/	??-???Q;�r&�@U�(3�+MS�K  �%q�+N6[!%i��%��?��%_EVN~ �4�-��6�2N

 }h3�UEV~ �!td:\ev�ent_user\�?B@C7GO/��YF|L:ASP@AEG�spotweldwM!C6�O}O�O*P�4!�?VO_I_�G �1_8_&_|_�_\_n_ �_�_o�_�_�_So�_ wo"o4ojo�o�o�o�o �o�o+O�o� 0��fx������zFWRK 2O��&!8�y��� g��������ӏ �.�	�R�d�?����� u���П������*��<��M�r����$V�ARS_CONFuI"�P
 FP�û���CMR�"2�V
�9��	�4ೠ��1: S�C130EF2 Q*���ę���x֊0�5��3�?��a0@a0pU0ȅ� )/h�r��ȓ�@��ҿ��Ϳ��k�O5�A���7ϲ�? B���R��� V�޿wϾ���jϿϪ� ��������=ߔ�� s�^�pߩ�\����ߓ��IA_WOQ�W<i��v,		�F�|(�6�G�P �I���H��RTWINU_RL ?&I����ߎ������������SIONTM;OUO � �B�XS۳�S���@�! FR�:\�\DATA��O  �� �MCA�LOGN� �  UD1A�E�Xr���' B@ �����`�����������x �� n6  �������6��  =���M�J ���g�TRAINМ�\�Bd�p�MQ����ңY&K (�ѝ	����� %[Im���������_GuE)�Z&K�`
���
� 
�?"'��R�E,�[�)����LE�X $\���1-e���VMPHASE'  &E�N����RTD_FILT�ER 2]&K �1��_� ??$?6? H?Z?l?~?�?�?��/ �?�?�?OO*O<ONO�`OrO��SHIFTMENU 1^�/
 <��%���O����O�O_�O�O C__,_y_P_b_�_�_��_�_�_�_�_-oo�	LIVE/SN�A��%vsflsiv�.?o�� SETU��bbmenuxo}oo�o�o�#�E)�_k�HMO�)�`.�z��ZD�ta\/
�<��P��$WAITDINEND��!rvvOK  ꩑|�r�S��yTIM����|G}���0�������xRELE�!@�vvs�<�xq_ACTU`?�t�x_J� b���%�o@����RD�IS����vpV_oAXSR|�2cYy�w�D(|�Ӡ_IR 3 �&t� 7
ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚϸ�Ͼ�NXVRy!�d7~�$ZABCv�1eY{ ,� �2����Oq��VSPT f7}�r{�
�j�o���j��ߣ�B�DCSCHb{ g�d���IPRrhY�6�H�Z��l���MPCF_G 1i��05׫�q�MP�j�6 �p5�����<��0  �ܳ�L?y?O����  �����3\�K4��+�+�&�'���Dd�8C��z��?�?�ۄ�4 �{��&�8�"J�1V���z�?����������/�� ��d��ðX�D̿73����W���3� FX?�����@��~�����P�0���C�Ą�{ k�W_�CYLIND�!l й� ,(  *���Ӧ0��/�  =/ O/a.��/��/�/�/ �/!/??&?i/J?�/ �/�?g?�?�?�/�?�?�O��2md� ġ�7OGLj�pO[O��O��'O�O�ז�AA��wSPHERE 2n��>?_�? _P_7_t_�?�O�_�_ 8?�__e_o�_:o!o �_po�o�_�_�o+o�o �o�oYo6HZ��ZZކ �ʆ