��   v��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@ � &�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  w�aIRTs1�	o`'2 L1���L1��R�	 �,��?���a�1`�b�ba �����y`� ��o��
 ��'�/SOFTP�@/�GEN�1?CUR�RENT=>�A,18,1�o1C�U �o�o,95,�2W���� �	(k}5	p�(�:� L�^�i��q9_��� ��Ϗ�����/��A�S�e���E,381��ğ֟�o� a��%�7�I�[�m� ��������ǯٯ�z� �!�3�E�W�i����������ÿտ���~a�TPTX��p���/�` s����$/soft�part/gen�link?hel�p=/md/tpmenu.dg�� �ϨϺ��υ����� &�8�J���n߀ߒߤ� ����W������"�4� F�X���|�����������a�f8�b�b�� ($p�-�@���T�?�x���a��a��c���c���� l���c��ah�ah�h�2�h�P.h��������q�`���`  ���|f ep��*h#h�Fd��g�Xc�B 1)hR �\ _� �REG VE�D]���who�lemod.ht}m�	singl	�doub �trip8browsQ��� ��u���//�@/���dev�.sl�/3� 1�,	t�/_�/;/i/ ??/?�/S?e?w?�?�?�?� H`�?�?  OO$O6OHOZOlO~O �F2P�?�O�O�O�O�O _�E�	�?�?;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo M'�o�o�o�o�o�o +=Oas�� �������?>� P�b�t���������Ώ ���O�����L�^� _'_�������ş� ����6�1�C�U�~� y�����Ư��ӯ�o� ��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�-��ϬϾ� ��������*�<�7� `�r�A�Sߨߺ�q��� i�����!�J�E�W� i����������� ��"��/���O�I�w� �������������� +=Oas�� �����,> Pbt���߼� ��//�����^/ Y/k/}/�/�/�/�/�/ �/�/?6?1?C?U?~? y?�?Y��?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ �R_d_v_�_�_�_�_ �_�_�_�o*o�_o�`oro�j�$UI_�TOPMENU �1K`�a?R 
d�a*Q�)*defau�lt5_]*level0 * [�	 �o�0��o'rtpio[�23]�8tpst[1[x)w9�o�	�=h58E01_l.png�~�6menu5�y�p�13�z��z	�14���q��]��� ������̏ޏ)Rr����+�=�O�a���p�rim=�pag�e,1422,1 h�����şן���@�1�C�U�g���|�class,5p�@����ɯۯ�����13��*�<�N�`�r���|�53������Pҿ�����|�8�� 1�C�U�g�y����ϯ� ��������"Y�`�a �o/��m!ηq�Y�w��avtyl}Tfqmf�[0nl�	��c[g164[w��59[x �qG���/��29�� o�%�1���{��m�� !�����0�B���f� x���������O�����@,>����2P �����\�� '9K����@��������1��@/$/6/H/Z/��|�?ainedi'ߑ/�/�/�/�/��co�nfig=sin�gle&|�wintp���/$?6?H?Z? !Z�a�h?�?�e�?� ;��?�?�?OO+O=O OO�?[O�O�O�O�O�O �O�O_a�%_L_^_p_ �_�_�_���_�_�_ o o$o�_HoZolo~o�o �o1o�o�o�o�o  2�oVhz��� ?���
��.�� @�d�v���������M� ����*�<�ˏ`�@r���������^� �;�M�sc�_;���As��X�}���e�u�� 0���P��t��h4�j�X�6e�u7�� ���ｿϿ���P� )�;�M�_�qσ�ϧπ�����������"�1�M�_�q߃ߕ� �Ϲ���������� 7�I�[�m����� ���������!�����6(�]�o��������$��74�������)t<ϯ\�5	TP?TX[209©|Dw24§J����w18�����02��A#��[�tv`�RdvL�0�K1���5S:��$treevie�w3��3��&du�al=o'81,26,4�O/a/s/ 2�/�/�/�/�/�/�/�?'?9?K?]?o?��;/��53$/6$���? �?�?
?#O5OGOYOkO }OO�O�O�O�O�O�OH�?�?��1�?6$2�8f_x_�_ �6_��edit��>_P_�_ �_o��/���_�So oo�o�oB�o�o��o A�o�+=O as��o���� ���(�9���Q�x� ��������ҏ�O��� �,�>�P�ߏt����� ����Ο]�����(� :�L�^�ퟂ������� ʯܯk� ��$�6�H� Z��l�������ƿؿ �y�� �2�D�V�h� ���Ϟϰ������ϕo �o��o@ߧE�c�u� �ߙ߽߬�����O��� �)�<�M�_�q��� W���������&�8� ��\�n���������E� ������"4��X j|����S� �0B�fx ����O��/ /,/>/P/�t/�/�/ �/�/�/]/�/??(? :?L?��߂?1ߦ?� ���?�?�?�?O$O5O GO�?SO}O�O�O�O�O �O�O�O��2_D_V_h_ z_�_�_�/�_�_�_�_ 
oo�_@oRodovo�o �o)o�o�o�o�o *�oN`r��� 7�����&�� J�\�n���������E� ڏ����"�4�ÏX� j�|�������a?s?� �?�sO_/�A�S�e� w������������� ��,�=�O�a�#_�� ����ο��=��(� :�L�^�pς�Ϧϸ� ������ ߏ�$�6�H� Z�l�~�ߐߴ����� ������2�D�V�h� z������������ 
����@�R�d�v��� ��)����������ƚԔ*defa�ult%��*level8�ٯw����? tp�st[1]�	�y��tpio[23���u����J\menu7�_l.png_&|13��5�{4�y4�u6��� //'/9/K/]/���/ �/�/�/�/�/j/�/?�#?5?G?Y?k?�"p�rim=|pag?e,74,1p?�?��?�?�?�?�"�6class,13�?�*O<ONO`OrOOB5�xO�O�O�O�O�O�# L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]o�oo�o`�$UI_�USERVIEW� 1֑֑�R 
��EDIT,Weld DATA ��double�����obmedit�1�o0BT�j�695�Pa�� ��m ��$�6�����cSTATUS�,POS�ftrip�o�o�o����ʏ܏��y2��+�=�O�a��33�_���� ��ϟz�ܟ� ���� E�W�i�{���0���ï կ������/�A�S� e��r������ѿ� ���ϼ�=�O�a�s� �ϗ�:ϻ�������� ���"�4ߦ�o߁ߓ� �߷�Z��������#� ��G�Y�k�}��:�D� ����2�����1�C� U���y���������d� ����	-��:L ^�������� );M_� ����v��� n7/I/[/m//"/�/ �/�/�/�/�/?!?3? E?W?/?v?�?�/�? �?�?�?OO�?AOSO eOwO�O,O�O�O�O�O �O�?__&_�Oa_s_ �_�_�_L_�_�_�_o o'o�_Ko]ooo�o�o 6b