��   ^��A��*SYST�EM*��V9.1�0214 8/�21/2020 A %  �����(�AMON_�DO_T   �$PORT�_TYPE  �@NUMJ/S�GNL7 L�$MIN_RA�NGI$MAX6rNOo ALxp �V�~ �COUN}TJ��AWE0�8 � $A�W0ENBJ $��G1LY_TI�V$WRN_A;LM�STP�
��E�C�.�W�TC�
J�AFT�_CHGxAVRG_INT��{�SAVE�YP~1ER_REG��T$WA� SIG6� OP��_VOLTS�����AMP�&A�E �#E_VL � &D'>% I*f$� �_ANL�  p 
$US0 S_CMD � �PRIORITY��"UPPER� �$LOW�$�#$�FDBK�"�RA�v �!SQ_AVG��#�#SD_� CE� � ��$ �܌ � LIN�!$�ARC_ENAB�L�!� 0DETE�C�!< ELD_S�P�$PD_UNI8��!92DIS�"��ID IM�#�1�  v1WFt2����CF�" � �$PS_MAN�UF �2O�DEL�5PROC�ESN0�0WFEE�W0ESC�2�2_F�I#1�1�1�7T _A�O�"�2I�6D�7D�C1�6L �"{2 ι CNV� 7 ?  $EQ�z,xODOU��2?@�TBd  �$?C 2 ��?@DD   �, � MM�!�$D� ��!?2 $F� �B֋4NV7	JBSE�L10_NOJDA�TA_s@�@ �{"WPpG
{M
��DWP7 �L@�L
 �WI�R_CLP4 �L@ASBU8  �H $4���R�4�YPRE�F� �U;A_ECU��  JB~ �S   $BP�EEPf#}!SCH>7 � �!���`�1e#dPK�*jFREQ.gULSwbSP�0fg2@y�!hyb*g�F�1;AI6 �ZCo VG}�hp dD�e�e�`P�	�a��dBVB�a�ZEROy}uS�LO]R�`NT�!P��cO	U\93�L FO7RMA0NAra�0�J3	� D�c�QWUXWSCCC @P8JU\�uT�IOEX7d� �A�Wfxcc�pS_91INp�� :1�UJ�� FAU�G"t0LO�0I�PD�!_�G]��R��A�p���STIC�@J�R�OBOT�ADY�H�ERRO�SE�d��`S�g�STA3RTE��!TR�0F~��CHDOG_�@�t��0_ACTIVtW��IH�TOR `OCOLL@�ӃC�0�1Q�2H��qE�2� ?Q:2TA�B�0 =�f5)$g1��RE��@92�I� �1R��r�%;E7��S�!S�UC*�N3FAILf��DSt@��LT��sABXP��NRDh2N3Px��RS�0�Y� N3�Q#�+3����)D�)D�)D���S�T�`3�3�3NO� ��B���Y�̤�0���R[2����� 91G�.�*�.��<�^� ;���-���.�S?�0��0PA� h������/HOUR_P��o � ��SE�0 �T<�:1HEpP6��GA�HPZ5�Y7�QLENGTH�"� `�P�#�����S�
BETO)F�0#SɦDn�w�x�.�UNy���91���2}!L�8  � �0���B���@������BISPp0E�RIC@�A)$F�SB� ��CURR �Bm4�!�dbg.���������0
`U!R�E}pd0W0������ NEW��2�PPIP�1_P9Oa�EK_Ӏ_R>��E_DBG`���Tp���3��4��5_QޕsEOTF7 � $��P�$�`x*�nfpNCi ?�cJ�f?�*dJ�*g ?�7fJ�7i?�FdJ�Fg0��Td��TfUP��9 ��qEPCR7A�� ��ل� L�Hr  ��%�4��00��2�X��0À3KIPTHE�RJ�ـ���KEf��0�&��WV�2��Eð;0�0��PHK-1��@��� RM��CH�S�PTL�0�$H�z�SW��BBONLC�$B��2pfbgF"WF �1t��q�zE"�!� s_W;6�AND1o�\�!ND2v3v�aS� �A� ����M~�� | $�0 �@g�e�*f�7b��Ff�TfADAP�!�LG�CSENS�Y�r ��EVP�!�� 4?p�Oֱ o3�$F�r�r7cr Fa�Tarm�'��&�{�&�!4�&5�&6�"��f��ʿܼ�� ��B��6B�6��46 ��65đ͒0�7w�����Pe@�V���TAI����)�A3T��	TX1�'EP>���\GP�0S��$��\O OVӀI��"[�AM!ܒK5M� AF��^1BEF֦LNd]�����%@��� mq `�ePPW)��:3�6i r��TRK�:�1�9MANU�qZ2m�D@DβOSR�EA � 	�y�&�`��  Ր�7y�q1^0Y6>H^1MIDU��If�!�����`�+�DEQ�w�CD0�!je�O �>P 4 ^'�q l&�S�������Q!�&P $ $E�LE�caQ�q5Ԇt	S_T�C����<;��r:�{:�0�TVPK �P� UU�uR�:�MU �eY�U��T� ���S$��S6XS��R���W������FW8�dBd��LAR�*�e *�)eO$`�O$p�O$��ЁQ_7�gUSh���cEC������PW{���_Og�#�e �f �eu)f��bw|�t���DI$�d�@Ewr~pLEw@|SIZ5RxVu�D��BOAR�C@h� ��� `��a p��r{a�r�Q�U$VENDր���OEVIC1xD D�#j~�JւV}�IN�`�t�1��q;�MA0�CwpFIB�URf�f�~,E p $,B�/�,B/2��F,�O���,BC��Ǳ��TO�ԩ�_R.@M�����މ$BUP�� 4 Аo�-����p��?!L��!�PU�RA�PREFLO]W�OSTi�Rwp�+���A�0�������&��S_DlqdM�ఽ�T��d'���MF ST/@���n��t M�A�Ԡf��ر�$���΂qADJD��#NE�Xc���4���T_P�!h��1M�b�#( �Æ8�S_!���$�HaO�!�,�PFL� GAP�2I� �����BJWT`�C�Y�p�x���[�!�s df�.s !r�@�-TOT�@�U��!U�IApT�WAR�~0V���Ahz��r�Y^v��<�KG?r��0��k��"XsNp  � 
PSCFl�"/( ��O���#�^��cQc�?!*�W�GLOBЯ"���� �NOT�!$��IXC9!�!AV��Y��\�$"�5�1p��W�_SHF[W$1X#Ɛ"I-�\� ?�t�RY�3`���p�3P��L@M�t���E�F UIFo�0�O|p��!�AD��\�APC�OUP����# @0��(�-�
 5�x��EQ{��@MMY ��T���T���
P�0�USTOz�� � ��{P}�� w
� �EMG� n�A% ,QMG��,� ��NOѠR�֨��7�����& !����э����s �Z2T�IR2T�qR��E�p�X`M���?�MI�T�CTSK�_WAIII��V�G	� S����7���T�_BUF����g�C`�ABNe��`��� ���������D>�=����GcSIN���R�E���1CT��NX���L�p�7���SsAVH��_PD��4I�e�W� LTn����PIP�s�0BG a`��[џ�fџ�qџ�v�P ��SPC�'� ,>#���b��Aҕ���� ���PP@A`z�����i2P��>�cHE�@i�?! k!k�r��bk�" j���"`�B��� SpB�R�B������_FIL�W�pB�UN�〷�b��F_@��.<�0wp��N�PSVO �C�0a��;PR>DIO�И�`s�p��TMB�^
PAP��� �󞢁_DYNe1i�W�r�F�`KEYe0G0��`@8�BF�1�@���� $#�RPR�O�U,$C"� �B@bCCAL��@`�`T��4i�P�_#!RTy#H���0A�� �$$�CLASS  /����! � � � � <0S�A�'�  ��!IRTU�0�/� �AWAO���A 4�!� � �!�!;EAɐ 2�(054;52�!?�Q338b51:5J5 J6�?�?�?�?�?�?�?�OO,O;96EXE <
01?C?U?g?y?�O �O�O�O
__._@_R_�d_?OɐS R!> gA�%�_�_�_�_�_o o'o9oKo]ooo�o�o��o��3NLG �2"< �q_qC?�lK<�!A��	mI	�; Bд!J X�5� 2�%��c�Gene�ral Purp�ose� MI�G (VoltsK, t�)�p\ ���p
AWMGEN�L.VR�vA*?EGLMG1�x�C1
�rBnu�Pxv�g �q�!�}<�N�`�r����sF�o�hCNV 2�	"<�2����sG 4� ��$����W�6�{��� l���ß�����؟� /��S�e������z� ��ѯ������+�=� �a�sL�=�����C� ܿ�Ϳ�$��H�Z� 9�~ϐ�oϴ��ϝ��� �ϣ� �2��V�h�G� ��k�}��ߡ�����w� ���@�R���v��g� ������������� 	�N�%�;���_�u��� ��������&J \;���gq�� ���F%V |[������ //�B/T/3/x/�/ i/�/�/�/�/�/�/? ,?��J?t?�/�?�? �?�?�?�?OO�?:O LO+OpO�OY?�O�O_O �O�O�O_$__H_'_�9_~_]_�_�_bNV�WP 2&��\�dT 
�_oo0o�d}USTOM 2}&�l  ;oP�o�o�o|	�d�e�nrDEFSVpR&���P<�o�s�Default SchA*w N`������ �+���a�s�J�y�𩏀����RFBKL�OG1 @[mTlaBG�����#��5�;�ۈ2���C�  s���������ۄ�LG_CNT  �[moa�RIOEoX 2[lDEe�A Ec��	�@=i�@=��Q
Wel?d Spee�a�c?IPM  �f� x���������ү����Eb $?���none=k�#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� ������������Rn� 2�\
�9��616-AU�G-23 13:�24:48�A�230816Ee�1324�C����Q)	Unde�finO�����
F�0��^����;��A>�#Wkm����� %	LA�BL�D_2=k@Ed�ac^��ig���āC 5��f���=h���19:�0����19C�C��D������� >�?�Wjd1C '�K���7/�U/c/�/��k`��/�//>��2D��3Eb̐m>?��.��V����/3T��
�_�1�? /�/{/A/�?OO6OzZNiAB���)37-ZO�O�/��?�� ��;?M?_?���O�?� x_�?AO;OO�_�_�_ �_�/�>oPo�L_o�Czo�o+)�o�o�o�o jon�>?Qcu �������� ��o�o>��o_���R� ��*����%� 7�I�[�m��������8ǟٟ�����C��OTF 2T�?����:�Տ^�p�G�ޝ==���*@��󭯿�I�PCR k2�paBH���*B��n��C����!�ffA� a =�+�OB�PMܠT�"�(R��W�uOܠT�#����������A��A��2345678901��퀠p_5�G�Y���à����@��,@�{���C��_h����S��SRAMOP 2���Q$������Y�RGS�EL R��   	Pr?ocess �?1��+ʼV�3�T�4
�9t�5�9h�7��F*��7�9���G0����ܠT�� ��"A|���A@�Z��B�&��Qh���Voltag�	ev�s�6<�DwF�X�@]yl�h���Wire feed sp����IPM�8<�� M�<�� �.�	�<�� ��*�<�N�`�r��� ��������������D��(R�z  �#��E�B��Q��o�����ݵt��V�����ѓCu�rrent�	Amp�u�<��? Q-?Qcu� ������// gh!��h%h!��h!�� h!��h!�h!�,�/ qװ��������!���! ���!���!��l/8}��?�����!Z�� )h/�	K/�?��?�?�?�?
��S R&�$��4ᨵ!O3OEM�?�:EO�O�O SOeOwO�O�O�O�O�O ;_M___+_�_�_a_ s_�_�_o�_�_�_Io [oo'o9o�o�o�o�o �o�o!�o�o'i {5G����� ��/����w��� ������я����� +��9M�k�a�k�}����)�ß�����������,9բUPܠ �୔=�o?��33:�>7�=L�S�>;���!��"���#��$��f�X'�$K��?^��>��r�� ?J2`�WIR/E 2!�<�������>�3�>��G(=�J*]�S?CFG "��v�@�#��|�������O����#�OUPLҠ#
���j������� w>��w;ۿO������ѿR�I�[̇�NB � Ƶ�� �UST_OM $�
6�c�ɿ �EMGOF�F %�6�#�LO*�&�ϑN��A�P�BM�� �uf�x  ���
,<�������ā�f���PCRg ' �~�@�bD�CE�5������D� _%��M�5p���%��