��   F�A��*SYST�EM*��V9.1�0214 8/�21/2020 A 
  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT  &F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBA�N��GI�eE�NC/  ~CRYPTE�  UOP��$$CL(   O���[!��	��u	P V� IONX(�  �}�l!IRTUA� �Z/�$DCS_C�OD?���_%�/  W�'_� �/��(S  �*�� $� 6�A91�"�!�	 $ b!��0=<?R?`?v?�? �?�?�?�?�?�?OO�*O8ONO\OrO��3S+UP� :�tO�O3F�O�O�O��  %\"Q���6_ �� V�[t&��j��T�O�_��LWJ_��� �V�_�KLUG�H 1�) � 9o)o;o Mo_oqo�o�o�o�o�o �o�o7o/AS ew������ ��+�=�O�a�s� ��������͏ߏ� � �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ���
�
�1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� "�7�I�[�m���� ������������3� E�W�i�{��������� ������,�AS ew������ �5