��  	G��A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ����AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO"  � A�LM�"ENB���&ON�!� MDG�/ 0 $DEBUG1A�"d
�$3AO� ."��!�_IF� � 
$ENABL@QC#� P dC#U5K�!MA�B �"��
� OG�f 0COURR_D1P $Q3GLIN@S1I4$C$�AUSOd�APPINFOEQ/� �L A �?1�5/ H ��79EQUIP� 2�0NAM�� ��2_OVR��$VERSI� �UP�0COU�PLE,   �$�!PPV1CESH C G1�!�PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1d��D�!U4 Q ��ARG1R�
 � $TIT1 d ��� 7Td7T� 7TTP7T55V65V75V85V95W05W>W�A�7URWQ7UfW1pW1
zW1�W1�W 6P!�SBN_CF�!-�0$!J� ; |
2�1_CMNT�$FLAGS]n�CHE"$Nbo_OPT�2��(�CELLSETU�P  `�0HYO�0 PRZ1%{c�MACRO�bREPR�hD0D+t@�تb{�eHM MN�B
1�UTOB� U�0 }9DEVIC4STI�0�� P@13��`BQdf"VAL��#ISP_UNI�#p_DOv7IyFR_F�@K%D13��;A�c�C_WAx?t�a�zOFF_@]N�DEL�xLF0pq�A�qr?q��p�C?�`�A�E��C#�s�ATB�t�d��WELDH2/0 =s�q"Q7ING�0$�QAx7PD2�4%$ASd3��BEl�P�_��BU�CC_AS�BFA�IL��DSB��F3AL0��ABN@��NRDY���`��zv��YN��SCH���pDE���yp���p�����|�STK>�0��	���	�NOj�?�ڂL��d�U* G��� 9 ���������߇ƗpƗ��ԘS_Fә1E��F�ƗSSŘ���P�1 �ON�F�HkOU�D�MI�1D�SEC`B�yi �HEK0~��GGAP������I� Ν GTH���0D_ȡ����T= ��륌� 
��p}�9!K���9!ƗUN14��5��#�MO� �sE �� [M�s��t�R�EV�B����QXiI� g�R�` � sOD}`��i�`M�m� ����/�"��� ŵ�!�X�@Dd p =E RD_E���?$FSSB�&W`kKB!�E2uAG� �J��  "��S�� V��t:5`�QCe`�a_�EDu � � C2�f�S�pa�l ��t$OP�@QB��q��_OK"�آTP_C� ���da�U �`LACm�^��J�<� FqCOMM� K�D��р@�p���OR��`BIGALLO�W� (K\��@VARw�d!�AB ��BL[@S � !,KJq��H`S�pZ@�M_O]�՗��CFd X�0G�R@��M�NF#LI���;@Uɠ�884�"� SWI�&"AX_No`����9���G� �0WARNMxp�d4�%`�L�Tb;�� CORz-rFLTRY�/TRAT T�`� �$ACC@�TB�� ��r$ORIأ.&�RT�`_S�FgϰCHGV0I����T��PA�I*��T���K�� � �#@a"�N�HDRՃ7�2�B�J; �CO�I�3J�4�J�5J�6J�7J�8�J�9�! Ȱx@�2w @� TRQ���$%f������_�U����e`COc <� ����
�3��2��LLEC��>o�MULTIV4�"�fѱA
2FS�IL�D���c� 
�1b w 4� STY2�bv�=��)2_��8C��� |9$�.pڰx�I`�* ��TOF �sE�	EXT3ء�B3�2�2�0���@�	1b.'.���
���  �"��/% �a�g�?s}@��A!��;AآM܁`Q  �TR>E� " L�0��	�`��pA�$J�OB��E����%IG� # d�,/>/ P(���#��B�_MORc$ t2�F͠�CNG�AŠTBA �6c�: /�9��0�19@G;aP/pH5�?�%L�����Bq�1��&rJ���_R������;J(@��8�<J� D81�@�9Q��2�@����}Rd&� 
�	�rG�R�`HwANC?$LGw� �a2q�͠���/���
0�2�R��Li�0�D��)�CDB`�C3RA�c�CAZ�`�H�ELT��FCT<�.�F"�`�)M#@�AI([O(X� ���
1�Rw�w 3�/�S���1��5�MP������HK&AEGS_SH�Q�W�ЅN0S��������'/  v@I#�Aq��Rc(��STD_�C�t�Q�3�UST��U��)kTITh�a~Ф	%�1IOy���@_Up�q��*c \����UpORzs `b��}�~p�`O~@N�SYR�G`�q�eUp��Љ�� ��DB�PXWORK��+�$SK��<����DB�TR�p , ��0A���c�B̎�W�DJDS _C`dд�sDPwPLzq �ё�s��DM�<wBY����2��H�9N�6p� q0DB�A��-�bHaPRi�M�
p��� ��. q�v�1$�$Z���L�y/��������0����P�� 1��tEN9E��� 2���~pREv��r3H� $C��.$L`�/$�s���tw�gINEV�a_D}�m�RO3���I;��~!�`�:���RET�URN���MMR�j"U琋�CʠNE�WMA`#�SIGN2��AJ@#�LA<�!��&P0$Po g1$P�@�24�M�;�O��S���a��o��v�Q�V�GO_AWT #�`�@`ъQe�`C)�o�CY� 	4'"�1�(����Ĕ2��2̖Na���C��4��DEVI�� 5 P $��RBU��PI̗P<��3�I_BY�;��J�T�1�HNDG�q6 Hv�c&�E�g㸣�#�㗣͖Џ`���`��L�70w��`�Ѭ�FBڬ(�FE�����͔��@�
ܱ8� �МQY�@�MCS4�Ƞ�dH���
�RHPWF��5:��J n����SLAVv.�9�INP���J��Ш����:P +B�S6@`�� �B�� 1�FI(b���	��5OaQ'OaW�	�NTV�V���SKI�CTE�*�@��b�]�QJ_�S�R_���SAF�v�5���_SV2EOXCLUv`-�%D~`L���Y��{�HI_VRP�RPPLY4px���u�۶���_ML�v`$�VRFY_s��M��IOC\�%C_�>PS�T�]�O/���LQSр��nt4Fqy�͓� �`P�en⯐6K�AUNF�����͕���ZqCHD`�$������ AF� CPU#��TFq��Wѝ_ס ;4��`T8��c�� aű9N�� <��8@�TЀ5� ��g�óSkGN=�0
$U0 ������Б� *0e �b��b��ANNUN�����͕U0�4v`'�w ����>P����LI�EF�`I�>���$F��&d`0OT��nt��prTq��lkq�`EM��NI�r!?'"|�G~�Aޱ���DAYecLOAD��ctu�os5kq�EFF_AXIɢ%@4�Yq�SO�����`_RTRQ�A� Dy�Q� Qt` E���� �@���WP  ���MuPC@E�� B��XT]2Xl�8FDUt�8E��bCAB��C8�*�NSj0ID�!WRBU�A:P�V%�V_T  �@��DI%0cD� �1$V�SE�T �2]3�1�o�
��]2f�1E_��lVEP	0SWAQ�0�� 3  A_0��O�HqPPAmI	RAa]2B�`�n�� ���S��@�@�%�� C�� ���RQDW�MS��P%AXt/lLIFEp�. uq:"�NA!^2J%��?#^2C�����C�P��N0�$ǁ�&��OV��V&sHE��]2SUP�!��:"p_�$��y!�_:3�%���'Z�*W��*�Q�'S�ሢ�RX�Z�@�q^1Y2=8C"��T�`��	N?�*��J%Q �_�@xH�I@�TE `��CACHt��3SCIZp&� ��%�NZ�oUFFI� � p��ct��os6kqx�M�P%DF 8��K�EYIMAG�TM���C#A��F��Ɓ���/�VIEK�aG��R�@LCĐ� �?�� 	I�?P�4H 6b�STo�!�B�Ѐ�DTp�D��D��@EMAIL�𽀣��^��FAUL�rI�R8���cPCOU�Pǀ�e,�DTO��QJ�< $�C5�S�T � IT��BUF@�7 ��7
�4`*`� 	B*T5�C�����BAcPSAVuU7R \2 :�U�W����P|T5�R�L��_*P[U5��Y#OT���`��P2�\p�Z?��WAXec+�=бX*P�éS_GA#
�� YN_���K E<� D0�!p���UM�� T��Fƀ�$݀��DI �E��`O�P��aL����GKQF�&�㌁�ax�����	�M�\��a�C&�SC_��K���`���d��RA�e�H�agDSP3F�bPC*{IM�S!sGq��a� �U�g� ��"��@IP`D��c{0 tTH[0���r��T��!sHS�csBSCQ�j0*�Vְ�z�p!c�tf���NV��G ��t[0v*PFAB`ds}`a�ǁSC�&��cME�R��bqFBCMP����`ET�� N6BFU� DUP���22��CDy�p�P6�C �ЀNO�х�O �������)PN�Cj�υR��@b�A���P��PH *ρL۰��� �QL����o�B���@� j�@���@���@��1@�7=�8=�9=�A ?��I�1V�1c�1p�1�}�1��1��1��1J��2��2I�V�2c�U2p�2}�2��2��U2��2��3��3I��3V�c�3p�3}�3���3��3��3��4����AEXT���Q Tb��Y`m&Y`:�d`����"�FDR�RT
PV���R:"�ɱ�r:"REM#F�U�OVM�c�A���TROV��DTl�P�MX'�IN��8� ��IND6�!
bȎ`B`W`G*a��!��@J%0D!�R�IV�n"GEA-R�aIO'K�lN}`����%(L�?@� >mZ_MCM50:!� �F� UR{�S� ,́MQ? ́ \p?4�@?4�Et�<ёgQX�R��T�0�Pa� �RI��I�7SETUP2_ U ��F6STD�px5TT���LѢלչ�7RBAC�NbV T��7R�d)§j%<��x`�IF�I�x`X�)�A ��PyTM�AFLUI~D�W �� `H PUR�`Q�"�R�a�p-PT�$ Iܴ$p�S$��?x|�J�`CO��P�SVRTl�G�x�$SHO#���CA�SS�p�Qp%�p��BG_���V���c���xp���}�FORC�B�,-�DATA��X��BFU�1�b"�2��a��/�[0��Y |�r�NAV`��p����S�Bn#�$VISI��vbS�CdSEZм�V*��O���B�IἉ ��$POt�I���FMR2>��Z Ȳ�� yɱ�`��ͷ������P��@�_���Ύ$IT_ᛄ"M��Ʋ���DGCLFރDGDY�LDDLѐ�5R&��J%W���~E[G@;	 T��FS�PD\ P�z��cB`$EX_.1`��"j3P5P�G�q���] �L�x�SW�^UO�DEBUG����GR��4@Un?�BKUJ�O1�7 O PO �мj���M��LOYOc�SMK E�R��AT�� _E ^� 7@��,�TE�RM %_)&�0OR�I�a% `)%��SM_�`��% a)%���h(bB)UPUBcg� -S��^p��7#� _��G�*� E�LTO�A�b�FIG�2�aЛ܀N$��$`$UFR�b�$À�!0��V OT7�TA�pɰ13wNST�`PAT�q<�0G2PTHJn����E�@�R���"ART��P�%�@�Q�B�aREyL�:9aSHFT�r(�aM1{8_��Rw���Jf& q $�'�0bvpʰ��\s9bSHI�0�sU9� �QAYLOvp2aHa1�]в�M18B�ׅ�pERVH�A f��8l�-7�`�2���sE��RC\�ׅA�SYM{aׅ�aWJ�'l�h�El�w1�If���U�D�`Ha{5� gF5PZs5@
��6OR�`M��Tw!��d��L001a�sHO���e �S1X��OC�!�>�$OP���a�.���䱩��d䰚PR�9aOU�sM3eV�RK5�U�X|�1��e$PWR��3IM�UIBR_�Sp40r�g `3�aUDlӳ3�SV	�eQ�df���$H�e!f`ADDR��H!GO2ata�ma��R���g Hz�SE���壬e�ec��ep�SE?��~��HS����h $gЈP_Dq�����b�PRM_R�|!H�TTP_H�i; (��OBJ��mb6��$��LE>3cP|)q�j � |�.b�AB_c�T#{rqSYP�s@�KRLi?HITCOU�t�� �P��P{r��l��P��PSSg�;�JQ�UERY_FLA��!b�B_WEBS;OC���HW���!��k�`�@INCPUdr�O:��qH��Q��dR��dR�p� ��IOLN��l 8�z�R��d�$SL���$INPUTM_!$�P��P��w ,}�SLA� m����مՄ��C���B�aIOpF�_AS�n��$!L��Ow���1��"b��!I������@HY���X�1�n��UOP�o `�v���F� H�F�O����PP&c�P�����O�ǒ���au�M��A6�p lH CTiA0BVpA��TI��`�E&P ��0PS�BU IDC �r���?��P>�|!�:�?0�qЂ��+����N��� ���IRCA|ڰ�� r �mymԀCY�`EA@��͡��ҬF�&c�k�R�g0�AA��ADAY_<G�B�NTVAE�V��.�Ȃk5:�.�SCA�*@.�CL��G����G���6�sr���l2����N_�PC⫠G��7�tЂ�Sޱ���JrG�>�p"�� 2s ���6��u���Jr�LABp?13� 9�UNI�9'�Q ITY���$xe�R���vЂM��R_URLT��$AL��EN�n�s�tg �Tv�T_Uk�� �J9�6�w X �����E��9�R����"] A�Ӂ��Jv���#FL9k���
Ӻ�
�UJR��x �mpFA�7��7<ҽD{�$J7�`O^�B$J8g�7PH!�p҂�78�c�8���f�APHI� Q�qӶ�D+J7J8�����L_KEd� � �Kt�LM��� y <��X�R�G���WATCH_VA��5@~�Fv_FIELDhey��L�ҁ�z R 51V>@¦K�CT��W�
�r�:�LG��{�� !��LG_SIZut���� �����FD��I������ ��" ���S����  ������" ��A8�� ��_CM#3`���g�-F�An�����r�T(���2�ိ�� ��������I��������" ����RyS�\0  (�SLN[р|���p �@ڂ��,��s:rYPLC9DAU_�EApt�|Tuk GqH}R�a �BOO�a?}� C7� `�IT�s�03�RE��SCR��s8��DI2�S0RGI"$D���+��TH�t �S[s�W�� �N+�JGMTMgNCH� �FN��bWK}��{UF���0�FWD�HL.�STP�V�Q X�� �RS�HP�(�C�4��B+�=P0T)Uq�/��>�a�@��Gm�0PO��'���i�sOC�EX'�TUI{I��ĳɠ��4	1�E3yd��0G���	�c���0�NO6AcNA ��QD�AI9�8ttt��EDCS��c��3�c�2O�8O�7S���2�8S�8IGN��G���zm��43DEOa5$LL�A{�HAT��~F�u�T��$��l�B�ä���-A\aF��P��PM�p�� 1�E2�E�3�Av��!�0 �m{Qk3������?�=Q�u� ����FST��Rv Ys�R0P� $E$VC $[[�p3VFV ��$ L4�F��P[�`=�[����Q$eENp�$d%6�_ � p- p`�� �S� �MC-� =�9�CLDP����TRQLI]���	i�TFLGR�P�a+cbr�D:�+g%�LD+ed+eORG��/!>b~U�RESERVU���d�c�d�b��S�c� � 	e/%dF+eSV 	`�	na��d�fRCLMC��d�o�oyw��a�M�p��Ѕ��$DEBUGMASI���	�Q�uTu05�E���TQ�MFR�Q��� � ~��HRS_RU����Q�A�T%FR3EQ��Q$%0��OVER-���o��F�A�P�EFIN�!%�Q�]qޑ�s�dǇ \���q��$9U�@޲?�`G�SPS�@��	�sC~ ��c�W�sU��bq�?( 	v�MIS�C.Ո d6�AR5Q��	��TBN�c ��&1ˈAX�R���·�EXCESH�ºQ��M���щm�a���T�R��SC�@� � H۱_�����S�����`J;PT�ċ &�i�FI��MI��� � �Po�]^H RCT�Ns�ȖOҚAҚ��Ԑ�C��u�ԐUSED�w O�@TЏ�PX ����������^P)�/��+eR� �pSZ��B�_FR�`T��\�Z_��^�CO>� P
HqK�čA�h�cu�B_��LICTB�� QUIRE=#MEO��O��)�1�L�PM�Ŏ �P���hr⛣�b��NDK����Џ4+��9�D�x�GINA�DRCSM\�S��0ё��S#��'�PSTLn�ѐ 4��LO̐f�DRI��EEX���ANGk2k��QOD-A�u���5�=���MFm����v�I�R�A�U&�( avSUP��U��F �RIGG>� � ��`�S '���SG&�T��R n�P~�P��r��#mqPGW�TI/�t᫐(�M\�Qr� t�MD��I)�ƕ0��q�Hϰk��DIyA���ANSW"P�mA�!�D})Hq�OR�b�`�Д 
��U��VB��`ײ2��O_Lp�ѕ �`�@�C��Np+����B��P�� ����P���KEI"��-$B8�p��zPND2r�a��2_TX�TXGTRA�31�%r���LOw ���$�G�T�,F�.�|�g�_�RR2����� .W�[A�a ?d$CALIĀ(��G�1��2�@RINܟ��<$R��SWq0t��%sABC���D_Jഡk���_�J3�
�1SPH��r�k�P�-�3,�(��vPk�\�J%sl�4�b�aO.AIM%p��CSKPj��> qs��J~��Q������8����İ_AZ�bh����ELAg�qOC�MPҳ�aJ���RT�q)Y�1�i�G�Ȁ�1�K40Y
ZWScMG ��3tJG�P�SCL���SPH�_�0����`k����RTER����S0��_�0�Q�A0S���DI��23U��DF^Pv�LWVEL	a�IN�R0&_BL �0k�.��l�J3<LDMECHPB%rF��IN� �q���|�H��2k� �sP_�� ����1��b?������DH�t3഑�v@$V��R��41$v �q�rV��$�a�Ro�����H �$B�EL �w�_ACCE4(�S'%qa ʐ)_� ����TJ��C-*�EX�RL6��& c�w'��w'.�W)�'�m#�'36�RO
�_��A!"� 1�uu�W!_MG�sDD!1��rFW�`��]#=5m#X"�28DE[;PPABmN�'RO� EE2 �A�?	`��AOqO�X!�^P�_��bSP.�pCTR�4Y}03 Z�a yQYN��A���6����1Mwq�ѭr�0O ��CINC a�̱Z2A4˂:G��́ENC� L��k��!XX"Ʉ+�IN�BI6���E���NTEN�T23_�r�CL!O�r�@�pI�U� �Fj��\��@ia�yC��FMOSI&1�y���1�s��PER�CH  k�q�  .Wұ9S���B3t��$��5)���A�"�UL �4��t����EF��J�V��FTRK��AY [�(�O��Q�"ecͰp/S�HB�pMOMcҀ˂O��`��T�Y3��0c�#�2��DU��7��S_BCKLSH_C�"�ewpV�p�3�j��caB�jA��CLALM�D}q>`��e�CHK�����GLRTY���ӁD��?�r��_�T_UMps�=vCps/1�Us�pLMT)�_L nt+�ywEs}�p�{rp�% �u�(>�aA�P�trXPC?QrXHI�۠%5�=uCMC7�/037C�N_��N6�4�t�S	FE!cYV�2��wG�p	��"x��CATD~SHþ�34iF?�xa�xFX�7�X�L "0PALDt8B_PCu'c_���� f"P��c&�uJ�A�T�a��?�'��TORQU�0/� Si�i0��R�i0��_W Ve�TU"!��#��#���I��I��I#F�尜�s�����+0VC"W 0�1Wd�1%�#089���+�JRK%�j�,]�u�DB� M��uНMP�_DL!�RGRV����#��#���H_^㈣� תCO1S�1 �LNl�� (�� 	�v 	�ۑE��3�����Z�V��M�Y����������T�HET0�ENK2a3#β#�CBӶkCB#C��AS�����۔�#�ӶSB8#$�޵GTS��1C0� �O�_Z�B�$DUp�W£�(5��DQnQ_�sjA+NE���!K$t;	��±AƵ����֥��LPH��§E��S(�@�3�@�B�� Q�j�T�q���V�V�� )�V8�VE�V�S�Va�Vo�V}�V��H�*�0�(ݭ�G�E�HS�Ha�Ho�H�}�H��O�O�OT��'�O8�OE�OS�UOa�Oo�O}�Oq��F���O�3�T��S�PBALANCE�_���LE;�H_ƵSP�$���3���>B�PFULC�������B��1�=U�TO_puT1T2	S"2N�a^"�@ 3�7a����"N#Ra�T�PO� `!��IN�SEG^"�AREV8X�@�ADIF�U��1���1��PO!B��a��dg2u��@�q��LCHWARL}2�2AB��feo��@��
AqXsX
aP�t)��� � 
p*��L!yEROB"P�CR�"l�� �C�J!_�T � �x $WEIGH@i@$ӥ)��IA�@IF�1;0LAG�2�rS�2� �27BIL�OD@`�@&�STd �P��`B� 1 �������
]@J"�1�  2y��D�DEBU��L� "~�MMY�9�%� N��m$i@3$D�!IQ$W $����  �D�O_� A�� <@�'& ���1��B��N�C�(_�@�0#�O�` �� E%\pT�@�A[qT�<O$� TICK�� �T1� %3�`(0N"P �#"PR�`�1��:5�F5� PROM�PCE� $IRk��1p�2�P�2�MAI��2A	B�5_���3� a@Rn��COD,#FU�0�ID_AP�5� {2~��G_SUFFېG ��1�152�DO=7x >5�=6GR��D[3&D�1E@�=Ev�D�$6 ���H� _FI+!9n�CORD� ��_"36�r�B�1� $ZDT�5� �%ߢ4 *�L_�NA�!(0�B:5DEF_I�H�B`6TF5 �96$962SF5@U`6IS��l��!��94yS"F3T�]$4=��rB"D �b�T,#Dh��O��"LOCKE ��C:?L?^7{QB@UME�BD2SD@U D�R&Bc%ES&DPT &B&{f{Q1C� �1E �B1E2S1C�g�eH� �P� iT� uQ��� Wh�X�e�S�TE�a��$� �LOOMB_r/w0�wVIS��ITY��A$�O�A_FR1IWs� SIuQYqB��R%0�w00�w3E#
�W\xWh{��^vn�9_�y;AEAS�;B@5�Vtŀ�P�2�v4~y�5~y6�ORMU�LA_I���G��G� h S.7�e%COEFF_O 1o r�1C�G���S�~"CA���/�#�!GR�� � �� $�PF�"X� TM�W܄�U2�S,���#ER� T�T�Dn6 �  ��LL<D:�PS�_SV�TH�$v6 �� G�6 �� ΂SETUuSMEA�0�0���!�B�� � q�] g @��������Q���B(0�Q�Q	�T���qFB�f1��P�Q�P����� N�0REC�A���!�SK_��� �P�1_USER�/�N�? s�N�/VEL�N�? v�j���I�@� �MT�!C�FGD��  �*0� ONOREȓ� ���� ��� 4 ���XYZ�C�@ J#��ʠ_ERR�� ����!�0���2!�:���� BUFIGNDX�Ȣ�pR7� H�CU��!�_��1�A����A'$Lt�OQ�軁@ ��GĂ� � $SI;��p�0�{R�VO�����PO�BJE����ADJ1U�"´ѰAY�AɳD��OU�@�_�\�1�B=^�Ta p.�v�-ǡ"DIR2��:�� ��ziDYNH�ry�v�T ��R^q�� ����OPWO}R�� �,� �SYSBU���SCOP��4�_���U��b� P�P����PAQ�������OP/@U�����)"f!�IMAG$��&�"3IMw�@�IN�p�~?�RGOVRDk���R��P�>�i� P�`�S��L�PB�|� ��PMC_E�@4�[!N��M��f!_"11d"� k�SL��E��� ��OVSL:�S�bDEX�QNP" �2g ��_k�� a@l��a@"�7�2�_"W�CZ�@�f�4�l�/_ZER���҃��D�� @נ��3O&�0RI±D
��0@�����ǡ�ܰLD��Z�T ATU9S��u!C_TV�C��B����Ṕ�Se!8���@E�� D�!� ��s�v3�A?�$���XE���\�p�;�b�㲠��UP��PoQPX�0.��]$y3��7��PG��}���$SUB���3]a����JMPW�AIT��'�LO�W�1���CVF�1+0RK���&�CCi�Rm�2_I�GNR_PL��D�BTB PsQB�W�0U��U� TI�G�j0ITNL�NS�R���R]pN<j0��PEED��	�HADOW ���ʰE����PS�PDD�� L�A`'�P"�0UN����.��Rw�q�LY(�@�  ���P��D���$���f0� 3LE��� PA�P����yP�~�>S�ARSIZ�4�@��CMQܰO>@�9�A�TT���-����M�EM�"f!�TUX���}��APL�0���� $���aSWIT�CH	�!WͰASr��1"LLB~��� $BAr+�D�S�BAM��h[Å)��w J5�䗡�"6�&Y!_KN�OW��"k�U�A�Dz(��-DQ��)PAYLOA���`3�_D�7��7Z3L�]aA��>PLCL_� !}�D2�!���Q4��_6Fi9C��?:��B4[�I?8R��?70�[4B�p�JLq��1_JI1i���AND/�
��4I2]1���qPLh AL_ �= -���!�Ѫ<pC�D3E��sJ3�0F� TU��PDCK��rR�C}O��_ALPH C�fCBE��(� O2L������� � ��� ?D_1:224D��ARc��H�Ex�F�C��TIA4Yu5Y6�MOMq�@S:S'S:S4S��B% �ADS^V'S^V4SPUB��R?T�U'S�U�4R���@G@�� � �M,2�� �1!A��� e$PIm���C@Z�7i`�'9iIkIkI+c�T�\f��\f����\Bg�Wª��HIGL#�& �f&\ K��f�c�h�\�i\&SAMP k�d�t�gs&� �3 o�Fq��z� Ut��_v�@ny�@z������P]u�q�b]uIN�|�p�c�x�{�t&�z�x�t�{�GAM�M�uS
���$G#ETW�@���D�D��M
��IB���I�$HI�_[�D�z���E����A������LW��̆Ì������ЩB�f� AC�CH�Kyг�ڐUNI_ �`����B�H�q�uY��RS��|VX�GC {�$BH 1���}I��RCH_DX�0����G��LEv�Z�в�嘩H���� MS�WFLV�QSCR&��10���SN�Wr3��:�|w�PnyN��]�PI3A�VMETHO}モ���+AX��h�X� ��N�ERI��t3C�IRB�5	�a�@F4�$q\s��ks��qLĐq�OOP\qp��0�kq��APP���F�И4�U�@��sRTբ�O�0�`��a����T`1����T`஺+`��)�MGڞ�,&SV~��PD�G� ���GRO<� ��S_SA�!��,ū�NO�@C��� �D�b��O?%?1h��o�W`�"_e���CDOA_�� UvP��u�h ��g��h����H3� >A0 M�U� 7� ^�YLc�1
�w��S�2Q��bׂ(����1��nӽ1_rđC�Z�M_WA�B�� �w����Mj  ��d0��A3)�	�(����PM��R� �� $Y�m��W"�n�԰L!51"��D  �D �D �4D{ ��AN� d�C#���pXj	O�C�qZ���P0 �TW� ���M��W� T�f�xϊϜ�P��ّ�,#�A_��� | SA���:Yl�'Sl�4S �Z����-ZR!\�*!(c!P���* 60P��P��PMON_�QUp � 8��QCOU���`Q�TH� HO[� H�YS�ES�" U�E µO5$� � ? P �|�3�RU�N_TO��A�O��b�P� P� `Cx��/���INDE��ROGRA��' o�}2��NE_NO��`IT�Q� D IN;FO��� ?!�
��m��@�OI��{ (p�SLEQ�f`��e� �. OS2�޻� 4�EN�ABN�^ PTIOyN���ERVEdbp[rac 3GCF<� @ J�Уqh+�h�R�\n���PEDIT��˓ �/��K�Q�c���E��NU��A�UT.��COPY��Q�`,ra:�M��Nx +*�PRUT�Ru "N�OUC�a�$Gep$��RGwADJ��� hS@X_��I͓���&��
�&W�(P�(�&�c� �N�0_CYCzN�pRGNS89�P��`LGO7�s@�NYQ_FREQ�RW�p�f-1SIZK8�LA��$1�!5S�p�eCREo���8��IFa�NA q�%k4_G��STA�TUS�VMAI�LrbA�1�LA�ST�1aA�$ELE�M<� �9�FFEASII�KrD� t��2���F٢�pn�I� l�$2�a���&KBAB2�@E� �`9V�1cFBAS�BdE�n��QU�`�`'�Y${A�GRM�PREC �qؐ�C���`��1�Dc � 2�S�[��	"B 2�  �s���tV�BW�B����p�ѡB3W�WߔDO!U�ӔO��$Pݡ�@=�GRID�2oBARS�gTYJΆ"OTO����� Q_�4!� �RnT�O��9� � ����POR��S��.�SSRV�0)�T�VDI0�T_e``#dPr`-g`-g4+i5+i�6+i7+i8a��F�?�<�O $VA�LU~C�D@pF>8�� !E;�ġ�S�1�۠AN�õb�1y�12ATO�TAL_�4I@rP�W3IvQ(tREG#EN&z;r��X�Hu0����f��TR�C�2�&q_S��w;pأV �!��rsdBE�3ݠ�B`��cV_HƗPDA��p�pS_�Y6���>6S�AR���2� h"IG�_SE�p�R�5_�d �tC_�V$CMXJ�C�T�DEE��
b�I:�ZS�-�N1�b�ENHANC'� p�AG�2A3��qINT`�!��F<Z��MASKʣ�@OVR����ݠ��1���WV��ayU��A�_'Fd{�V�PS�LG%��a� \ ��?57��p�0S8���4f�Us�V�|��s��7aUP�TE|���@� (cq⟦J3�.�N3IL_�MM4�VQB۠��T!Q�𖣷�@C����5V�C-�P_�'��7�MN�V1M�V1�[�2j�2[�3j�3
[�4j�4[�����ޣ��ޣ����IN��V�IB�'�����2��2#�3�3#�4�4#���6�O�2����D`�Q`����P�L�0TOR ��I�NƵ��R��L���T $MC_F,  5���L ����pM?�I���OS� ]��f���KE�EP_HNADD" �!B�h@L�C�ᐐAbĮQ�t�c�O��A� ���pcë�c�REMz�bĺ1�R��Զ���U�4eb�HP�WD  B�S�BMӁ�PCOLL�AB���`e�qq2�� IT0��&"NO�FCALE����7� ,��FLK��A�$SYN��`�M���C@���pUP_�DLY���ODE�LA�л1�2Y��A�D��  �QSK;IP$�� ��Pb aOp਒(���P_b  ��ד ��� �׵ � s �D`��Q`��^`��@k`��x`�څ`��9�!O�J2R� ���AX�@T'3���A���� >¡�>���RD�C�aT�� ��R�˸R`1ɺȲ
T�RGE�4CгXRFcLG���ŐSWX�
TSPC��!UM�_��ؓ2TH2N�RQk�� 1ݏ 	���Q8 � D� ��:�l@O2_PC�#��S��|�A.0L10_CL2q���́ ��  b�'`����F(������� ��+U��г +� �b9�lCHЅ�������~DESI�G��'UVL1��1���Hs10��_DYS�(�����F  ;11�� l3�i�0��o�F&�AT��q$ ]Q07�'+$�  �����HOME(� �2����p��! �3��DVhz�V� �4���`���	// ��
�5��>/P/b/t/(�/�/-'6��/�/0�/�/?? U�!7��8?J?\?n?�?�?-'8��?�?�?��?�?O-%S���  �A�Pp6�����E�T� T0���D	v�CIOՑ�I�Ip@5�OB�_OP��ESr�C��POW=E��� �@_�r���"t �Z��BR$DSBf�GN�AOs��Cq�`�����Z�CIk _T_SPE%�z�CMD�W��Â�a��ޘ�DBG_\@PU������SEq�̀ �2�4C=��2S23�2�E� ���7E|o���ICEUSs<�U�ARIT�qq�OPB.ЭbFLOW�TR�@r���PƮaCUV` �aUX�Tҁ�a��ERFAiC;d��U�`-"wSCH��� t3�0���QH�@�$�p�pOM���A�  t���UPD����qPT�@Y�EX��x�c!�FA�e�G��r>fq � �цpZ�� (�AL� ��3u���:R;�  2�� �S���@��	� �$X���_�GROUQ�sT�\ ��vDSP�vJ/OGLI�cF����,a7�N�����ސ�f=K�`_MIR�q�Tf�MT��AP�`�c�*�Z�`�SYq��t�]��@�BRKH��avl�AXI~A  f�@�q��rρ�<�u�BSOC�v���N��DUMMY1�6,�$SV��D�EQnSFSPD_�OVR.����DL؂�sOR�P@N��b�Fv���pOV�u;SF�RUN����F8��a�sUFRAvN�TOldLCH�Ҍ���OVׄ8��pW�- ��sy�P�����_�8�� @E�TI�NVE$PKAOFS2ǐCSp��WD ���`�����R#�ÀTRO��R(�FD��(�M�B_C4��B� BL~���q0�6��qP�V�adB�` ���G1�D�AMB�$��`r�����_MH��b<��C���T$����q~CT�$HBK�a/�ءI�O_E�Q��PPA۪�������R��DVC_�PdCI�@q`RI�҆a`�1h���`�3h���"��`��pׁUdC�p�FCAB��^B[�"��&�k��h�O�UX/�SUOBCPU_R�pS�� ���Z��`��I�Z��?R��$HW_C@� t`���N��N@�pNp�$U-�z�|t�m�ATTRIEМ���pCYC��ұC�A���FLTR_2_FIqCsY��fVz��P�{CHK_�`�SCT�F_m�F1_w� ҉�FSeQR�r�CHA����A�Q�{b@�RSD��bQ��s`QP_To�? ��L�q`EM�@��Mn�T.��Np.��Ӷ��DIAGuRAI�LACV���MpL�O��f�<�$P�S�r`B �����P�RJ�SZ�& �Ct<�C 	��FUN��aRIN�Z�Y@0��?�����S_�pu àh�@Ѥh�-�Ѥ?CBLCUR}��aA������DAx�0i�����LD�`ˀ�����qr� ���T�I��}�Np$C�E_RIA��oRA�F�P�SG�[ L�T�2��Cs��C�OI<��DF_L�@P���as`LM�SF;H�RDYO�ѐRG� �Hb��Y@����MULSE����Ǽ�.s�$J�J�����FAN_ALM�MWRN!HACRD`@�ffs�2�Vaz�R�_��/�AU�R�R3ԇbTO_SBRU��p�
m�>�|G�MPINF���������REGF`FNV�`�Sb�DP�N�FL_Ž�$�M�����c��Np�(/C�P� ��dA���PӐa��@$�qA$Y�R�a�}r�S�� ��7�EG&P�sˀ�A�P�D��25������D�AXE�wROBn�zRED�vWR�P2k�_���SYh��tϠ&S!'WRI�P�M�STOP�s�`l�J�Eo��@�6��Df�pBa ��h&7��.��OTO��@Y�ARY�s�"�ѝ��B��pFIM��s$LwINK��GTH�"M
pT_^#���98���!XYZ�b�*9�&OFFŐ�"�P�� �(� B�p4�`D4��mP�`E3FI���^7K�nSÄ4��t_J,aNr���#��[ w$�*30��9`Е1��2�2C#Q4�DU�³��3%���TUR X"�E�!�X0 `�7FL� l�̳�$@5�d)35�Ғ 1��@K�pM/��6��������cORQ@�ֺqn�8��J�O �N��E���q��DOVE�A�RM�`�Aj 
Up
Uv	VaWαWpTANE��!
Q L�Q�A�IP��QU��AW�Up�U.S�qE)R�qr�	 �E��Dp$��TAQNpa5`�`�ҫ'��׶��AX�� Nr�ᝰV��"+e��7i ��7i��6j�6jq 6j@� 6j� 6j06j1�0 6f��3i��Ci��Si�� ci��si���i��i���i��i�a�iDEBUE�$@�L��tqڒ�"AB��ء ��C9V͠D� 
�rq� r�u5��w���w���w ��wq!�w�!�w�!�w�1R��0L��"E3LA�B[2�EA�N�GR�O���2E��B_ �ѸVM$��U0� l���p�E��y��ANDr@� ��T���%�Qy�  ��M^ �������� �NT, ��+�VEL���eT5���=���E3NmAc�� �$���ASS  �������� �x�ʐSI����]��㆔�I��x������AAVM, �K 2 ��� 0  G�5������.%� %�	H�9�\�����J���n���8�����G�������АBSQ� 1���� <�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ���������������/�A�S�e��L�M�AX�� h��n5�  dz�IN�����y�PRE_EX�E������D���|��АIOCNV*B�� ȑ�P���0���1��IO_�� 1]ݛP $͠�r�0]��Z��?�h��� }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	���-�?�Q�c�z�LAR�MRECOV ������6LMD/G FQ k��LM_IF  F��h��"�4�F�T����wωϛϭϾ�, 
 ����b�n ��1�C�T�$��x� _ߜ�[�����������s�NGTOL  ��� 	 A �  >�P�z�PPI�NFO Ż� Ķ������  �»��者��� ��6� �2�l�V���z����������� (:L^p������غPPLIC�ATION ?�-�����ArcToo�l  
V9.10P/30O���
88340�-F0S@10�5-"47D�F1(�Non}e�FRA�� 6p�_A�CTIVEp�  ��7�  �UT/OMOD ��5���CHGAPON�L$/ 8#OUP�LED 1��� u y/�/�/�CUREQ 1	�W  T�)�,�,�	�/	5� 4����"_ARC �Wel��AW����"AWTOPKS6HKY?���/ �/�/?v?�?�?�?�? �?�? OOO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�o 0BTfx��� ������,�>� P�b�t���������Ώ ����(�:�L�^� p���ܟ����ʟ��  ��$�6�H�Z�l�~� د����Ư�����  �2�D�V�h�z�Կ�� ��¿����
��.� @�R�d�v��ϚϬϾ�0�����̹%TO(�/�#DO_CLEA�NE/�|�NM  -� �/������� ��.DSPDgRYR��V%HI" ��@��~������ ������� �2�D�V��MAX� c��1T't�Xc�sp"s�PLUGGc d�p#�%PRC5�B��"��m�_���O��>��SEGF< ^0 .7�߶�~���8���1LAP[�n 03 2DVhz��������T�OTAL����USWENU[ h+ I��M/2� RGDIS�PMMC^021C�+3�@@�"h$O�Y�{�I�RG_S�TRING 1
~4+
�M- �S�
�!_ITwEM1�&  n� �/??%?7?I?[?m? ?�?�?�?�?�?�?�?�O!O3OEOI/�O SIGNAL��%Tryou�t mode�%�Inp�@Simu�lated�!O�ut�LOVE�RRX� = 10�0�"In cy�cl�E�!Pro?g Abor�C�!��Dstatus��D�@cess F�ault\Ale�rT	Heart�beaSgCHand BrokeZE WOY_k_}_�_�_�_�_�_�__��+_��/ �_9oKo]ooo�o�o�o �o�o�o�o�o#5�GYk}�_WOR : �+�q)o���� �%�7�I�[�m���� ����Ǐُ����!�3�PO�+1QY��{ B�|�������ğ֟� ����0�B�T�f�x����������үT�DEV\���p��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h�>z�PALTm�� �{����������#� 5�G�Y�k�}ߏߡ߳������������GRIy��+E���m�� ������������� !�3�E�W�i�{�������3�+ Rm��]��� #5GYk}� �������1CU��PREG �Ύg���� �/!/3/E/W/i/{/ �/�/�/�/�/�/�/[M��$ARG_�pD ?	���<1��  �	$[F	[�P8]P7�[Gq9/0S�BN_CONFIQGj@<;�A�B�1��1CII_SAVE  [D�1�3/0�TCELLSET�UP <:%  OME_IO[M�[L%MOV_H8�0	OOREP��ZO�%:UTOBACK��1<9�2FRwA:\{ eO,{�0'`�@{�H�� �K�0 �23/08/�13 15:18:50{r8{_0-_Z_Q_�L��z_�_@�_�_�_�_�_{��_ )o;oMo_oqo�oo�o �o�o�o�o�o7 I[m��������!���� � �A_}C_\AT�BCKCTL.TMH�`�r�������oKINI���E�5�1~z@MESSAG�0�ρ�1D0ڋODE_QD�0�6�5�O����wCPAUSm� �!�<; ,,		�r0<5q��e� �������������� ��S�=�w�a�s������D�N�TSK � T��O��z@UP3DT�͇d���XWZD_ENB8̈́�:'�STA̅<1��.1WJ@ODP�2�<;4W��)13-AU�G-2P7:33 P42O��˿ݿ�1��F�L��߿*�7�`����
u�B��� ̐  :�f������j�ROBGR-PҨ�A�"��WEWELp�������6:56��D
/LAB_��_�D������9k�f��n� �߭���qσ���+47XIS�0UN��Ԧ��1��� 	 �I���Ck�`� 	1! ��pګ{ V��D�1�2��t��{�V�Q�� �AN� ��n�� �$�)�Z��������0�3�ME�T��2D鄰 P�U�@n��@ ��G@�6?�@�f@,�@vo���>��>����='�?3�^�>l�m?��&9�SCRDC�FG 1<5�A ���  ���);M�O{Q�9������ ��^�?Qc�u�� :'7}AG�R=��2��C�NA�#@;;	}D�_[EDˀ1�������%-I�EDT!-���m/���@!(~BI/:r2p_F�B/�/  ���%2 �/6K�/F?7��+?? �/�/n?�/�#3�?'? OK?]>�?KO�?�?:O�?�#4�O�?�OO]>��O_^OpO_�O�#5 O_�O�_�O]>x_�_*_<_�_`_�#6o�_ho �_]>Do�o�_o�o,o�#7�oWo4{o]>@{�o�oj�o�#8�[/ ��^=�G� ��6���#9��̏�^=���Z�l�����!CR�/"�� ��X}r�ݟ$�6�̟Z���% NO_DEL���GE_UNU�SE��IGAL�LOW 1���   (*S�YSTEM*L�	$SERV_���Lٗ�POSREGƠ�$£Lܗ�NU�MŪ�حPMU|C�L�LAYO��L�PMPA�LS��CYC10�$�7�!�%�]�UL�SU�٭9� ���Ls���BOXOR=IɥCUR_��ح�PMCNV����10M���T4�DLIB����	*�PROGRA��?PG_MI%�O�Fa�AL/�n�X�a��B�ϗ�$FLU?I_RESU=���ϯ����MR��������Wr?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7��I�[�6�LAL_OUT ���#�WD_ABOR>��g���ITR_RT/N  �Ā���?NONSTO ��� O�CE_RIgA_Id���0 �� FCFG �*0��9_P}A��GP 1CU���$��C;��� ��-C� C � (� M�+C8� @� H�  �CX� `� h� p�� x��� �� �
� �� �Rdv����?�HE�O�NFI����G_mP߰1C  1�����/ /2/D/�V/h/�KPAUSf��1��0 M� j/�/���/�/�/�/? �/6?H?.?l?R?|?�?@�?�?�?�?�?r,M��NFO 1���S  � 	p�OO;�=O ³����B������5�$��6���B��*��ƌA��u�K�zbC3��{\V�AB�3� �O=C�Ǹ�COLLECT_=�+F��R�GEN�/����R�ANDE��C�GR���1234567890[W:ұ�SY_kVF��
 %}�;�)�_ �_���_�_o���_�_ Too1oCo�ogoyo�o �o�o�o�o,�o	 t?Qc���� ����L��5V��;2�K ]9RIO !DYQ�ǁ��Ώ������TMRr 2"�� ��1
-���#��<���Y_MORz�$w ��ŕdAřݟ ˟��%����m{��%��,�?����x�;�K��;ѷ� R�=&�O������C4/  A����;�=�A{�Cz  B��$B�"  �@Ң��;�:dYڍ��ARI=S'���?�z�(���/�d���T_DEFz� �X�%J�������N�US<��0��KEY_TBL  ��06B�	
��� !"#$%�&'()*+,-�./dW:;<=>�?@ABCe�GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������h���͓���������������������������������耇����������������������}!b�LCKp��	b���STA�����_AUTO_D�O��&�IND8T��_T10�"׃T2o�V� T{RLd�LETE�����_SCREE�N �k�cscU MM�ENU 1)�� <o�|�D�UE#�M� ��i�k�������� ����6���l�C�U� ��y�����������  ��	V-?e�u ����
�� R);�_q�� ��/��<//%/ r/I/[/�/�/�/�/�/ �/�/&?�/?5?n?E? W?�?{?�?�?�?�?�? "O�?OXO/OAO�OeO wO�O�O�O�O_�O�O�B__�_MANU3AL���DBc�j������DBG_ER�RLj�*�D�C Q_�_�_n�Q�NUMLIM���[���
�QPXWO_RK 1+��_�_oqo�o�o�oS�DBwTB_�� ,�]�ģ����o�DB__AWAY�SD��GCP ��=��1b�b_AL`��bB�RY���ը��X_�PW 1-��h�
No`���|��f_MLГIS�
{@{��sOoNTIM��������vGy
��\sM?OTNEND��[t�RECORD 1�3� ����G�O���u���
r�� ŏ׏鏀�����<� ��`�r����1���)� ޟM���&�8�ӟ\� ˟�����ȯگI� ��m�"���F�X�j�|� 믠��Ŀ3����� ύ�Bϱ�M�տ�Ϝ� ����/���S���w�,� >�P�b��φ�q�߼� +������s�(��� ^��߂���=���� K� �o�$�6�H����� ~������������� �� ��D��hz����bTOLER7ENCtB�Qrp�L�͈PCSS_�CNSTCY 2�4?i��P�Or� 	);Q_q� ������//�)/7/I/[/�DEV�ICE 25� �f�/�/�/�/�/ ??,?>?P?b?���HNDGD 6���`Czu:O��L/S 27�-t?�? �?OO,O>OPOv?��PARAM 8�hy8rwUbD�5�5SL?AVE 9�=�7_CFG :�O�bCdMC:\�� L%04d.CSVaO"�c	_!�>�A 6SCH>P�1��bNI_~_�G�bF�nR�Q�_�Y�Q�@JCP��S�^"��a�>�_CRC_OUT� ;�-�afO_N�OCOD�@<hw~�MSGN =^��G�#M�1�3-AUG-23? 16:179P�A�vj5:199P�&? Wzz�i�a�bN�`ra�M��?Þ�j��a�n��CVERSION� ejV4�.2.11�{EF�LOGIC 1>^� 	�X�@�Iy�QY}+rPROG�_ENB<��6ysU�LS�w �6+r_�ACCLIM�v���C��sWRSTJNT�F��A�+qMO�|�QPb�tI?NIT ?�
^�v�A �vOPT�@� ?	6��
 ?	R575bCc��74h�6i�7i�50��t��2i��X��|%wF�TO  R���o�&vV�DEX��wd�riP$�PA�TH AejA�\�q����HCP�_CLNTID y?	v�C �[�Zß�IAG_G�RP 2D�I �> 	 �@K�@G��?���?l��>� �ٚ���8�ٜ5��� a�O�?ϧb�?> ��i��^?�Vm?S���ٙf403� 6789012�345����� ��s��@n���@i�#@d��/@_�w@Z~��@U/@O��@I��@D(��ٚѠiQ@�6TpX6P�� A�� � 9PB4ٜ� ٔR��iQ
Т1��-�@)hs@$���@ bN@���@ڠ��@?�D@+2�	���-�2�A�2�P�R���@N@I��@D�@>�y@9��@4���.v�@(��@"�\��������п�V�L�@Gl��@BJ@<z��@6ڠ0�`@*��$���@��&�8�J�\�V��=q@���F@|�@3�3@�R@-�?���?��`?�+�ϲ���������̑҂��-�@&�@�����!?�?� �,�>�P�b� t�V� �(�:��^�p� ��D��������x� ����6�H�&�l�~�� ��:���q�����Ѥ��x������Y�?��?�z���(�o5AF4� ��L4R� �(�@�p�8�Q��@-: I �m@����%�Ah.�=H��9=Ƨ�=�^�5=�v ��>��(�=�,v��,�^ �iQ�C)�<(�U�Rc 4�����ٙA@hR?0���"�� 0Vh4��t�8�����
/��>���y,"�R=�?��=��z<!(�o��G�T/G�(�@8U8U����(�$@9P���*��uB��J���B�B�?�B%�(��T$�/�.'�p5.�*11n,�\��=�-���c+�a Bk B��BC�A��@�Z?؟�?�iQ<�P��O�ոdֿx��83B��6����?�0��30��1C�;
���$��iPu� �?O O9O�(TOZB�ٙ�99�4�B�ܻ��$O �O O�O�O�O�O�O#_�2�>���>ˠ������>����@V�?j��_��'_u_�CT_�CONFIG �EDo�ceg��U�STBF_TTS�w
�y�S p�st��V5`MAU�p���rMSW_CF��PF��  )��jO�CVIEW�PG'm3���ןyo�o�o �o�o�oPrgo�o  2DV�oz��� ��c�
��.�@� R�d����������Џ �q���*�<�N�`� �������̟ޟ� ��&�8�J�\�n����������ȯگ�|\R%C cH`��R!���� $�Y�H�}�l�����ſ�dSBL_FAULT I�<h߱GPMSK�W�P�TDIAG J��Y�!�S��Q�UD1: 67�89012345 O¬RC��W��Pb_�� �ϯ���������	�� -�?�Q�c�u߇ߙ߫�j�?���
z��߂V�TRECP(�:�
 H�:�a���y�v��� �����������*� <�N�`�r��������������=gUMP_OPTION�P���TR b�S�P�ME�UY_TE�MP  È�+3BQ0m �L1W�UNI`�Um�Y�N_BRK K�Ro=fEDITOR���F�_�EN�T 1L� � ,&
LAB_WELD_�5մ1&��:ֲ�(e L�p����� // /=/$/a/s/Z/ �/~/�/�/�/�/�/? �/$?K?2?o?V?�?�? �?�?�?�?�?�?#O
O�GO.O� MGDI_�STA�+am�N�CsC1M'k �P���O�O��
��d�� _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o&�o �o�o�o�iQ�o" 4FXj|��� ������0�B� T�f�x��j�o����͏ ߏ�o��'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uϏ�}ϫϽ� �������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� �ϙϣ����}����� �!�3�E�W�i�{��� ������������ /ASe��� �����+= Oas����� ��//'/9/K/]/ o/��/�/�/�/��/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgO�/�O�O �O�O�/�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oyOko�o�o�o�O�O �o%7I[m ������� �!�3�E�W�qo�o�� ����Ï�o����� /�A�S�e�w������� ��џ�����+�=� O�ɏ{���������Տ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�s�}� �ϡϳ�ͯ������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�k�Y������ ��������)�;�M� _�q������������� ��%7Ic�u� ��Y����� !3EWi{� ������// //A/[mw/�/�/�/ ��/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKOe/ oO�O�O�O�/�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCo]Ogoyo�o�o �O�o�o�o�o	- ?Qcu���� �����)�;�Uo G�q������o�oˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�M�_�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+ϥ� W�a�sυϗϱ����� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�O�Y�k�}� ��ϳ���������� �1�C�U�g�y����� ����������	- G�5cu���� ���);M _q������ �//%/?Q[/m/ /5/��/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO 7/I/SOeOwO�O�/�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'oAOKo]o oo�o�O�o�o�o�o�o �o#5GYk} �������� �9oC�U�g�y��o�� ����ӏ���	��-� ?�Q�c�u��������� ϟ����1�#�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ��� �)�;�E�W�i�{ϕ� �ϱ����������� /�A�S�e�w߉ߛ߭� ����������3�=� O�a�s�ϗ����� ������'�9�K�]� o��������������� ��+�5GYk�� ������� 1CUgy�� �����	/#/ ?/Q/c/}s/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�?��?O/ �$EN�ETMODE 1�N~%� W + + &%�HOZK*@RROR_PROG %7J�%%&�O�IxETAB_LE  7K�/��O�O_WxBSEV�_NUM FB  �AA=PxA�_AUTO_EN�B  dE?CuD_;NORQ O7KYA}<R  *��P���P��P��PHP+��P�_�_�_nTFLT9RZ_lVHIS9S)!�?@g[_ALM 1]P7K �&$�\% +�_no�o�o�oȶo�o�__2RtP  �7K�QZBz*@T�CP_VER �!7J!�O�o$EX�TLOG_REQ�f�eY_sSIZ\hZtSTK�y�U��\rTOL  �)!Dzb�A= Zt_BWD�`�p��V�q_B�sDI�q ;Q~%�sXD<)!�{STEP��|*@0�OP_DO��(AFDR_GRP� 1R7I�Qd 	���Z@��n&����c?���$,MT�� ��$ ����ن�������Bt��B|�
B����Bu|�B
��FBA<`�AA��A�� Bc���B�HA5?�7A�Ԧ��� r�]���������ޟɟ�  @��As?�>(���+ 
 K�f�A�	��ћ��Eb؟�ҟw�b���*�@  ~��@�33@�Ǡ	ˣ�@¡毄������F@ 5�E���@�5�%��L��FZ!D�`��D�� BT���@����?� y ��#�6������5�Zf5�ES����(#� %"��YUV��XH��KFEATURE� S~%�p^A�ArcToo�l �)"En�glish Di�ctionary�*�4D Stan�dard#�Analog I/O"��A5�e Shif�tw�rc EQ �Program �Select��S?oftpar�ǝ��Weld��ced�ures���Co�re���Rampwing_�uto���wa�Updat�e(�matic ?Backup(�V��ground E�dit �-�Cam�erar�Fv�Ce�llr�{�nrRn�dIm[Ӓ�omm�on calibg UI����sh�������c�	���ne,�	�ty��s�����nt���Monit�or=�ntr�e�liab��)�DH�CP˒�ata ?Acquish��?iagnosR�o����ocument? Viewet���ua��heck ?Safety��-��han�� Rob��rv��q!���)ʊF�s��F���-�x�t weavS�c�h%�xt. DI�O��nfi"�|�e�nd.�Errs�L(���i�s��rm���� �p'�FCTN �Menu�����T�P In��fac\�-�Gen��l���Eq L��8ig�E'9m�p Ma�sk Exc*�g�r�HT% ��xy �Sv��igh-wSpe.�Ski��������mmuni�cQ�on��Hou�r ���s�(co�nnX�2�ncr' stru>��
!�e���J��-�KA�REL Cmd.� L� ua�XR�un-Tiq�EnQvN��:�+U�sS��S/W*�Lice�nse�����Bo�ok(Syste�m)'�MACRO�s,�/OffseZ�MMRm�i����MechStop"��t�����i����1&x.�o�S�D.od��wit��g(i���y.�ƅ+Optm�/�#��fil��'g���ulti-T�  �+�ORNTBASE Fun+>-�PCM f"8(��Po��� �I=Re�gi�r��,6ri0��!9~9p�Nu����<�8��Adju� �>x���=tatu}1��?��,�RDM0�o}t;�scoveD��)Eea� q�Fre�q Anly��Rem' ��nR�)E5B85�9�ues�ńG�o��r )�SNPX� b�#�SN% CCli���N��P rC�D�OU� 8$P�Eo�=t ssag յE���O!p 0��V^�/I&]UMILI�B�_`RP Fir�m9�p^PAcc<n�v�TPTX��^Teln��_aQ���q]or�@ SimGular��!fu��AP8�XZmЍ�#&��gev.]U1�ri���_USB po,����iP��a��f?R EVNT�o�`nexcept.�`j@W4�ej�P�VC��r��-(V��.r�_h?u�K9{S�@SC�U�qSGE�|uUI�&�W��8�|b PlF�~5���� (���������6�uZD?T Appl�'�x�f�s�Grid9Aplaym�mPZԇ�R%r.R�����F�< A�200i��c��larm Cau�se/h@edE�A�scii��Loa9d��1�UplG���yc��~�0�`� �RAe`���yQ�NR�TL�_4nline Hel��-6'�,6{0x1��tr"�6�4MB DRAM���FRO ������c� PB� .'�ma�i���K�RR�6L��Sup�b�!}9à��} croL4C�E��9vrt�4C&�� 3�*�<�i�`�r����� ÿ��̿����/�&� 8�e�\�nψϒϿ϶� ��������+�"�4�a� X�j߄ߎ߻߲����� ����'��0�]�T�f� ������������� #��,�Y�P�b�|��� ������������ (UL^x��� ����$Q HZt~���� ��// /M/D/V/ p/z/�/�/�/�/�/�/ ?
??I?@?R?l?v? �?�?�?�?�?�?OO OEO<ONOhOrO�O�O �O�O�O�O___A_ 8_J_d_n_�_�_�_�_ �_�_o�_o=o4oFo `ojo�o�o�o�o�o�o �o90B\f �������� �5�,�>�X�b����� ��ŏ��Ώ����1� (�:�T�^��������� ��ʟ��� �-�$�6� P�Z���~�������Ư ����)� �2�L�V� ��z�������¿�� ��%��.�H�R��v� �ϵϬϾ�������!� �*�D�N�{�r߄߱� �ߺ���������&� @�J�w�n����� ��������"�<�F� s�j�|����������� ��8Bof x������ 4>kbt� �����/// 0/:/g/^/p/�/�/�/ �/�/�/	? ??,?6? c?Z?l?�?�?�?�?�? �?O�?O(O2O_OVO hO�O�O�O�O�O�O_ �O
_$_._[_R_d_�_ �_�_�_�_�_�_�_o  o*oWoNo`o�o�o�o �o�o�o�o�o& SJ\����� �����"�O�F� X���|�������ď� �����K�B�T��� x������������� ��G�>�P�}�t��� ����������� C�:�L�y�p������� ���ܿ���?�6� H�u�l�~ϫϢϴ��� ������;�2�D�q� h�zߧߞ߰�������  �
�7�.�@�m�d�v� ������������� 3�*�<�i�`�r����� ����������/& 8e\n���� ����+"4a Xj������ ��'//0/]/T/f/ �/�/�/�/�/�/�/�/ #??,?Y?P?b?�?�?��?�?�?�?�?�5 � H541��3A2FR782� G50 EJ614�DG76 EAWSP�,G1[GRCRPH8�\FTUgFJ545�DH[FVCAM EC�LIO�FRI�GU�IF,F6�GCMSyC�HgFSTYLDG�2�FCNRE,F5�2[FR63+GSC�H EDOCVLVC�SU EORSFR�869DG0OG88�FEIO�FR54�7FR69[FESE�T�GrGJqIWMG��G�WMASK EP�RXYX7 FOC��F�P3�H7F�PCH3�fJ6BH53{VH�EhLCH�VOPLn�VJ50/fPS�gcMCfG�`�W55OF�MDSW�g"gOP�"gMPR�F<PSh0�CFORBS fCMb�G0w�POG50Sg[51�G51Ox0�F�PRS�W69fF{RD�FFREQ,F�MCNVmXH93�CFSNBA�GFgSHLBVM�w<P3W�NN_h2CFHTC�gFTMIV4@{VT{PA�FTPTX(�#EL�v�`{W86G4@�FJ95�FTUTv#g95fUEV�VwUEC�VUFR�F�VCCψOFVI�PVCSCW�CS�G'VaPI�hOFWE]BgFHTTgG62W�WIO�Ry�CGv:�IG�IPGv�IRCVDG"gH�75�FR66��7��WRMz2/fR]j4�f��OF�@FNVD��VD0��F�AL�O�VCTO�GNN�fM}xOLXENuD,FLڇFVR�E �8������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿���  OH541��2#�oR782$�50$�oJ614T�76$ɯAWSP4�1s�RkCRd�8t�TU���J545T�s�VC{AM$�CLIO�ʻRI��UIF4�6���CMSC4܃�S�TYLT�2��CN�RE4�52s�R6�33�SCH$�DO�CV��CSU$�O{RS��R869T��0c�88#�EIO�C�R54C�R69�s�ESET�˒�JΑ�WMG$��MA{SK$�PRXYd�M7$�OC�`�3��hC�`�S�3��J6R��53��H�LCH��OPL��J506��PSb�MC��p��c�55c�MDSW����OP��MPR�ڠ��0S�ORB-S��CM#�0`�c�50�51��5u1c0��PRSS�69��FRD��FwREQ4�MCNT����H93S�SNByA$��SHLBTڱM2�Г�NN#�2�S�HTC��TMI�c�@���TPAC�T7PTX�EL�
p����8B�@�#�J95n��TUT��95��wUEVS�UEC��wUFR��VCCc,�O��VIPc�CS�C�CSG����I�d�c�WEB��HTuT��6��WIO�*mR�CG�+IG�+wIPG#
IRCcڻDG��H75��R�66�;7B�Ra2
��R!�4��0c�0�n#�NVDS�D0�;�F!LALO��CT�O��NN��M�O]LR�END4�Lr+FVRC�ȺO�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�o 0BTfx��� ������,�>� P�b�t���������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l�~� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� ��������*�<�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�?O  O2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�� ��STD~�LANG(� #�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����'�9K]o��RB=T'�OPTN��p���
+DPN&�@"/4/F/X/j/|/�� �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h?z?  ��?�?�?�?��?�?�=99E��$FEAT_AD�D ?	����/A7@  	�8@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������������""DDEM�O S/I   �8i_q� �����
 -7d[m��� ���/�/)/3/ `/W/i/�/�/�/�/�/ �/?�/?%?/?\?S? e?�?�?�?�?�?�?�? �?O!O+OXOOOaO�O �O�O�O�O�O�O�O_ _'_T_K_]_�_�_�_ �_�_�_�_�_�_o#o PoGoYo�o}o�o�o�o �o�o�o�oLC U�y����� ����H�?�Q�~� u������������ ��D�;�M�z�q��� �������ݟ�	�� @�7�I�v�m������ ���ٯ���<�3� E�r�i�{�������޿ տ���8�/�A�n� e�wϤϛϭ������� ���4�+�=�j�a�s� �ߗߩ���������� 0�'�9�f�]�o��� ������������,�#� 5�b�Y�k��������� ��������(1^ Ug������ ��$-ZQc ��������  //)/V/M/_/�/�/ �/�/�/�/�/�/?? %?R?I?[?�??�?�? �?�?�?�?OO!ONO EOWO�O{O�O�O�O�O �O�O___J_A_S_ �_w_�_�_�_�_�_�_ oooFo=oOo|oso �o�o�o�o�o�o B9Kxo�� �������>� 5�G�t�k�}������� ͏׏����:�1�C� p�g�y�������ɟӟ  ���	�6�-�?�l�c� u�������ůϯ��� �2�)�;�h�_�q��� ������˿����.� %�7�d�[�mϚϑϣ� ����������*�!�3� `�W�iߖߍߟ߹��� ������&��/�\�S� e���������� ��"��+�X�O�a��� �������������� 'TK]��� �����# PGY�}��� ���///L/C/ U/�/y/�/�/�/�/�/ �/?	??H???Q?~? u?�?�?�?�?�?�?O OODO;OMOzOqO�O �O�O�O�O�O
___ @_7_I_v_m__�_�_ �_�_�_o�_o<o3o Eoroio{o�o�o�o�o �o�o8/An ew������ ��4�+�=�j�a�s� ����ď��͏���� 0�'�9�f�]�o����� ����ɟ�����,�#� 5�b�Y�k��������� ů����(��1�^� U�g������������ ���$��-�Z�Q�c� }χϴϫϽ�������  ��)�V�M�_�y߃� �ߧ߹��������� %�R�I�[�u���� ����������!�N� E�W�q�{��������� ����JAS mw������ F=Ois ������// /B/9/K/e/o/�/�/ �/�/�/�/?�/?>? 5?G?a?k?�?�?�?�? �?�?O�?O:O1OCO ]OgO�O�O�O�O�O�O  _�O	_6_-_?_Y_c_ �_�_�_�_�_�_�_�_ o2o)o;oUo_o�o�o �o�o�o�o�o�o. %7Q[��� �����*�!�M�  D�c�u� ��������Ϗ��� �)�;�M�_�q����� ����˟ݟ���%� 7�I�[�m�������� ǯٯ����!�3�E� W�i�{�������ÿտ �����/�A�S�e� wωϛϭϿ������� ��+�=�O�a�s߅� �ߩ߻��������� '�9�K�]�o���� �����������#�5� G�Y�k�}��������� ������1CU gy������ �	-?Qcu �������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� �������������'9K	   LQgy���� ���	-?Q cu������ �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?m??�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� ������� #5GYk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{������� ��������/A
PU Hk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/��A�S��$FEAT�_DEMOIN [ X�����X�}k�INDEXx�����k�ILEC�OMP T�;������f����SETUP2 �U��Â��  N �_A�P2BCK 1V~��  �)T�D"�1�%�U�X��� C���V����;�П_� ݟ���*���N�`�� �������I�ޯm�� ���8�ǯ\��i��� !���E�ڿ�{�ϟ� 4�F�տj����Ϡ�/� ��S���w���߭�B� ��f�x�ߜ�+����� a��߅��,��P��� t����9���]��� ���(���L�^���� �����G���k� �� 6��Z��~� �C��y�2 D�h���� Q�u
//�@/� d/v//�/)/�/�/_/ �/�/?�/%?N?ȉ���P � 2�*�.VRU?�?0*��?�?
3�?�?�%�0P�C�?#O0FR6�:OON�?sOKT ���O�O8E�O�Lz�dO<�O�&*.F�?*_"1	:C_W\�O{_
[STM�_�_7B=@D�_�]j_�_
[H�_�2o�W o�_�_�oZGIF�o�o�U�oaosoZJPG<�U`(�o�o�JJS�Ŀ0Rs�j%
�JavaScri3pt�CS�C���V0�� %Ca�scading �Style Sh�eetso�� 
A�RGNAME.D)T��<�P\��p���q�󏟏�DI'SP*��.ބ9����	�i�w�#�
TP�EINS.XML���Ώ:\��x�ځC�ustom To�olbar��*�PASSWORDn�~�.FRS:\>����_�Passwo�rd Config��/ȯW�����4? "���F�X��|���� ��A�ֿe�������0� ��T��Mϊ�Ϯ�=� ����s�ߗ�,�>��� b��φ��'߼�K��� o�����:���^�p� �ߔ�#����Y���}� ����H���l���e� ��1���U�������  ��DV��z	�- ?�c���.� R�v��;� �q/�*/��`/ ��//}/�/I/�/m/ ??�/8?�/\?n?�/ �?!?�?E?W?�?{?O �?	OFO�?jO�?�O�O /O�OSO�O�O�O_�O B_�O�Ox__�_+_�_ �_a_�_�_o,o�_Po �_to�oo�o9o�o]o oo�o(�o!^�o ���G�k � ��6��Z����� ���C����y���� 2�D�ӏh�������-� Q��u������@� ϟ9�v����)���Я _������*���N�ݯ r�����7�̿[�ſ ϑ�&ϵ�J�\�뿀� Ϥ϶�E���i��ύ����4���$FIL�E_DGBCK �1V��!���� < ��)
SUMMA�RY.DG>����MD:r߲����Diag Sum�mary����
C?ONSLOG�ߋ�����6���Con�sole log�7��	TPACC�N,��%y�����TP Accou�ntinX���F�R6:IPKDM�P.ZIP����
��;�����Exception?�����MEMCHECKЬ�����J�Me�mory Dat�a���!l�)	FTP)������L�mment� TBDG�L �>I)ETHERNET<�΁�����Ether�net N�fig�ura^���1DCSVRF;!3L���% ve�rify all�O�M.cDIFFD*<����%fdiff�����CHG01���V/a�~/�- )2L/3/E/ �/�{/�/"3�/�/�/^? �/�?6�VTRNDIAG.LS�?;?M?�?z���1 Ope�� Log ��no�stic�וɿ)VDEV�2D�AT�?�?�?�?b�VisADevisceOKIMG�2�1�AOSO�O�#~DI�mag�OKUP�/@ES.O�OFR�S:\._o]��U�pdates L�isto_���@FLEXEVEN���O�O�_a�Q UIF Evb	@�_�  ,�t)
�PSRBWLD.CMo��ZR6oq_�K�PS_ROBO�WELh�:GI�GE	Oo�_�o���GigEXo�NߵA�)�aHADOW�o�o�o|���Shadow Changes���a�<rRCMERRtYk �����pCFG Er�ror�@tail>� MA����pSGLIB���8��rI� St� A�-�>��)r�Z�D�o��o����Z�D@ad��3� <rNOTI��������Notif�ic�3�(f�AG ��������;��� _����$���H�ݯ �~����7�I�دm� ���� ���ǿV��z� �!ϰ�E�Կi�{�
� ��.�����d��ψ�� ��*�S���w�ߛ߭� <���`�����+�� O�a��߅���8�� ��n����'�9���]� �����"���F����� |���5��Bk�� ���T�x �C�gy� ,�P���/� ?/Q/�u//�/�/:/ �/^/�/?�/)?�/M? �/Z?�??�?6?�?�? l?O�?%O7O�?[O�? O�O O�ODO�OhO�O _�O3_�OW_i_�O�_ _�_�_R_�_v_oo �_Ao�_eo�_ro�o*o �oNo�o�o�o�o= O�os��8� \���'��K�� o������4�ɏۏj� ����#�5�ďY��}� �����B�ןf���� ��1���U�g������ ����P��t�	���� ?�ίc�򯇿��(��� L��󿂿Ϧ�;�M���$FILE_F�RSPRT  ���1�����\�MDON�LY 1Vp�(�� 
 �)M�D:_VDAEX?TP.ZZZN��������6%N�O Back f�ile ��(�S�6)ܿ7���[�$�h� ��ֿ��D�����z�� ��3�E���i��ߍ�� .���R���v������ A���e�w����*��� ��`�����+��O ��s��8�\ ��'�K]�����`�VIS�BCK��x���*�.VD�/pF�R:\�ION\�DATA\���pVision VD�./<v/�/ ��/��/_/�/?�/ *?�/N?`?�/�??�? 7?I?�?m?OO�?8O �?\O�?mO�O!O�OEO �O�O{O_�O4_�O�O j_�O�_�_[_�_S_�_ w_�_o�_Bo�_foxo o�o+o�oOoao�oV��LUI_CONF�IG Wp�|�{ $ �c��{p�Xj|����y@p|x�o�� � �2�B��e�w��� ����D�������� +�O�a�s������� @�͟ߟ���'��� K�]�o�������<�ɯ ۯ����#���G�Y� k�}�����8�ſ׿� ���϶�C�U�g�y� �ϝ�4���������	� ���?�Q�c�u߇�� �߽���������)� ;�M�_�q����� ���������%�7�I� [�m����������� ������!3EWi {������ �/ASe�v �����z// +/=/O/a/��/�/�/ �/�/�/v/??'?9? K?]?�/�?�?�?�?�? �?r?�?O#O5OGOYO �?}O�O�O�O�O�OnO �O__1_C_U_�Oy_ �_�_�_�_X_�_�_	o o-o?o�_couo�o�o �o�oTo�o�o) ;�o_q���� P����%�7�� [�m��������L�ُ ����!�3�ƏW�i��{�������A�͐x���ʓ�$FLUI�_DATA X�������D��RESU_LT 2Y��#�� �T�/�wizard/g�uided/st�eps/ExpertٟZ�l�~��������Ưد�������Continu�e with G7�ance�W�i� {�������ÿտ���,�� ˒-̑��><�0 �M�<������\��.�ps ϧϹ��������� %�7�I�[�m�,�M��� �߸������� ��$� 6�H�Z�l�~�\�N�`��r���torch ������*�<�N�`� r���������y����� &8J\n� ����������>��wproc��H Zl~����� ��/��2/D/V/h/ z/�/�/�/�/�/�/�/�
??��7?{����@�TimeUS/DST&?�?�?�? �?�?OO,O>OPObO~%�EnablE� �O�O�O�O�O�O__�&_8_J_\_n_˒�8�F?�_j?|?�624 �?�_o"o4oFoXojo |o�o�o�oqO�O�o�o 0BTfx� ���_�_�_�_w��-�?�Region �R�d�v����������Џ���!�America<@�R� d�v���������П����!��qy��P�8�$��2Edi��� ����ʯܯ� ��$��6�H�Z�+ Tou�ch Panel� �� (reco/mmen��)h��� ��ѿ�����+�=�O�a� ��0�B���f�|x��2acces/� ����/�A�S�e�w���ߛ߭�,Con�nect to Network�� ����)�;�M�_�q����$���p��ϚϬ��\!�ϐ0I�ntroduct >�Q�c�u��������� ������ /);M _q������� 0?��0 
��R#����� ��//(/:/L/^/ �/�/�/�/�/�/�/� ??$?6?H?Z?�x3P:H�?l�? �?�?OO+O=OOOaO sO�O�O�Oh/�O�O�O __'_9_K_]_o_�_ �_�_�_v?�?�?�_�? #o5oGoYoko}o�o�o �o�o�o�o�o�O1 CUgy���� ���	��_*��_N� ou���������Ϗ� ���)�;�M�_�p� ��������˟ݟ�� �%�7�I�[��|�>� ��b�ǯٯ����!� 3�E�W�i�{������� p�տ�����/�A� S�e�wωϛϭ�l��� ���ϴ���+�=�O�a� s߅ߗߩ߻������� �¿'�9�K�]�o�� �������������  ���D�V��}����� ����������1 CU�y���� ���	-?Q �Z�4�~�j��� �//)/;/M/_/q/ �/�/�/f�/�/�/? ?%?7?I?[?m??�? �?b���?�?�!O 3OEOWOiO{O�O�O�O �O�O�O�O�/_/_A_ S_e_w_�_�_�_�_�_ �_�_�?�?�?�?LoO so�o�o�o�o�o�o�o '9K
_o� �������� #�5�G�Y�o*o<o�� `oŏ׏�����1� C�U�g�y�����\�� ӟ���	��-�?�Q� c�u�������j�|��� 𯲏�)�;�M�_�q� ��������˿ݿ￮�  �%�7�I�[�m�ϑ� �ϵ��������ϼ�� �B��i�{ߍߟ߱� ����������/�A� S�d�w������� ������+�=�O�� p�2ߔ�V߻������� '9K]o� ��d����� #5GYk}�� `��������/1/ C/U/g/y/�/�/�/�/ �/�/�/�?-???Q? c?u?�?�?�?�?�?�? �?�O�8OJO?qO �O�O�O�O�O�O�O_ _%_7_I_?m__�_ �_�_�_�_�_�_o!o 3oEoONO(Oro�o^O �o�o�o�o/A Sew��Z_�� ����+�=�O�a� s�����Vo�ozoď� �o�'�9�K�]�o��� ������ɟ۟ퟬ� #�5�G�Y�k�}����� ��ůׯ鯨���̏ޏ @��g�y��������� ӿ���	��-�?��� c�uχϙϫϽ����� ����)�;�M��� 0���T���������� �%�7�I�[�m��� Pϵ����������!� 3�E�W�i�{�����^� p߂�����/A Sew����� ����+=Oa s������� ��/��6/��]/o/�/ �/�/�/�/�/�/�/? #?5?G?X/k?}?�?�? �?�?�?�?�?OO1O CO/dO&/�OJ/�O�O �O�O�O	__-_?_Q_ c_u_�_�_X?�_�_�_ �_oo)o;oMo_oqo �o�oTO�oxO�o�O�o %7I[m� ������_�!� 3�E�W�i�{������� ÏՏ珦o��o,�>� �e�w���������џ �����+�=��a� s���������ͯ߯� ��'�9���B��f� ��R���ɿۿ���� #�5�G�Y�k�}Ϗ�N� ������������1� C�U�g�yߋ�J���n� ���ߤ�	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������߮� ����4��[m� ������! 3��Wi{��� ����////A/  $�/H�/�/�/ �/�/??+?=?O?a? s?�?D�?�?�?�?�? OO'O9OKO]OoO�O �OR/d/v/�O�/�O_ #_5_G_Y_k_}_�_�_ �_�_�_�?�_oo1o CoUogoyo�o�o�o�o �o�o�O�O*�OQ cu������ ���)�;�L_�q� ��������ˏݏ�� �%�7��oX�|�> ����ǟٟ����!� 3�E�W�i�{���L��� ïկ�����/�A� S�e�w���H���l�ο ������+�=�O�a� sυϗϩϻ����Ϟ� ��'�9�K�]�o߁� �ߥ߷����ߚ��߾�  �2���Y�k�}��� ������������1� ��U�g�y��������� ������	-��6� �Z�F���� �);M_q �B������/ /%/7/I/[/m//> �b�/�/��/?!? 3?E?W?i?{?�?�?�? �?�?��?OO/OAO SOeOwO�O�O�O�O�O �/�/�/�/(_�/O_a_ s_�_�_�_�_�_�_�_ oo'o�?Ko]ooo�o �o�o�o�o�o�o�o #5�O__z<_� �������1� C�U�g�y�8o������ ӏ���	��-�?�Q� c�u���FXj̟� ���)�;�M�_�q� ��������˯��ܯ� �%�7�I�[�m���� ����ǿٿ������� ��E�W�i�{ύϟϱ� ����������/�@� S�e�w߉ߛ߭߿��� ������+��L�� p�2ϗ��������� ��'�9�K�]�o��� @ߥ����������� #5GYk}<� `�����1 CUgy���� ����	//-/?/Q/ c/u/�/�/�/�/�/� �/�?&?�M?_?q? �?�?�?�?�?�?�?O O%O�IO[OmOO�O �O�O�O�O�O�O_!_ �/*??N_x_:?�_�_ �_�_�_�_oo/oAo Soeowo6O�o�o�o�o �o�o+=Oa s2_|_V_���_� ��'�9�K�]�o��� ������ɏ�o���� #�5�G�Y�k�}����� ��ş������ C�U�g�y��������� ӯ���	��ڏ?�Q� c�u���������Ͽ� ���)�����n� 0��ϧϹ�������� �%�7�I�[�m�,��� �ߵ����������!� 3�E�W�i�{�:�L�^� ���������/�A� S�e�w���������~� ����+=Oa s�������� ����9K]o� �������/ #/4G/Y/k/}/�/�/ �/�/�/�/�/??� @?d?&�?�?�?�? �?�?�?	OO-O?OQO cOuO4/�O�O�O�O�O �O__)_;_M___q_ 0?�_T?�_x?z_�_o o%o7oIo[omoo�o �o�o�o�O�o�o! 3EWi{��� ��_��_���oA� S�e�w���������я ������o=�O�a� s���������͟ߟ� �����B�l�.� ������ɯۯ���� #�5�G�Y�k�*����� ��ſ׿�����1� C�U�g�&�p�J��Ͼ� ������	��-�?�Q� c�u߇ߙ߽߫�|��� ����)�;�M�_�q� �����xϊϜϮ� ���7�I�[�m���� �������������� 3EWi{��� ��������  �b$������ ��//+/=/O/a/  �/�/�/�/�/�/�/ ??'?9?K?]?o?. @R�?v�?�?�?O #O5OGOYOkO}O�O�O �Or/�O�O�O__1_ C_U_g_y_�_�_�_�_ �?�_�?o�?-o?oQo couo�o�o�o�o�o�o �o(o;M_q �������� ��_4��_X�o��� ����Ǐُ����!� 3�E�W�i�(������ ß՟�����/�A� S�e�$���H���l�n� �����+�=�O�a� s���������z�߿� ��'�9�K�]�oρ� �ϥϷ�v��Ϛ���� ҿ5�G�Y�k�}ߏߡ� �����������̿1� C�U�g�y������ ������	������6� `�"߇����������� ��);M_� ������� %7I[�d�>� ��t����/!/ 3/E/W/i/{/�/�/�/ p�/�/�/??/?A? S?e?w?�?�?�?l~ ��O�+O=OOOaO sO�O�O�O�O�O�O�O _�/'_9_K_]_o_�_ �_�_�_�_�_�_�_o �?�?�?VoO}o�o�o �o�o�o�o�o1 CU_y���� ���	��-�?�Q� c�"o4oFo��joϏ� ���)�;�M�_�q� ������f��ݟ�� �%�7�I�[�m���� ����t�֯������!� 3�E�W�i�{������� ÿտ�����/�A� S�e�wωϛϭϿ��� �����Ư(��L�� s߅ߗߩ߻������� ��'�9�K�]�ρ� ������������� #�5�G�Y��z�<ߞ� `�b�������1 CUgy���n� ���	-?Q cu���j���� �/�)/;/M/_/q/ �/�/�/�/�/�/�/? �%?7?I?[?m??�? �?�?�?�?�?�?�/ �*OTO/{O�O�O�O �O�O�O�O__/_A_ S_?w_�_�_�_�_�_ �_�_oo+o=oOoO XO2O|o�ohO�o�o�o '9K]o� ��d_����� #�5�G�Y�k�}����� `oro�o�o���o�1� C�U�g�y��������� ӟ�����-�?�Q� c�u���������ϯ� ��ď֏�J��q� ��������˿ݿ�� �%�7�I��m�ϑ� �ϵ����������!� 3�E�W��(�:���^� ����������/�A� S�e�w���ZϬ��� ������+�=�O�a� s�������h������� ��'9K]o� ������� #5GYk}�� �������/�� @/g/y/�/�/�/�/ �/�/�/	??-???Q? u?�?�?�?�?�?�? �?OO)O;OMO/nO 0/�OT/VO�O�O�O_ _%_7_I_[_m__�_ �_b?�_�_�_�_o!o 3oEoWoio{o�o�o^O �o�O�o�o�_/A Sew����� ���_�+�=�O�a� s���������͏ߏ� �o�o�o�H�
o��� ������ɟ۟���� #�5�G��k�}����� ��ůׯ�����1� C��L�&�p���\��� ӿ���	��-�?�Q� c�uχϙ�X������� ����)�;�M�_�q� �ߕ�T�f�x����߮� �%�7�I�[�m��� �����������!� 3�E�W�i�{������� ��������������>  �ew����� ��+=��a s������� //'/9/K/
. �/R�/�/�/�/�/? #?5?G?Y?k?}?�?N �?�?�?�?�?OO1O COUOgOyO�O�O\/�O �/�O�/	__-_?_Q_ c_u_�_�_�_�_�_�_ �__o)o;oMo_oqo �o�o�o�o�o�o�o�O �O4�O[m� �������!� 3�E�oi�{������� ÏՏ�����/�A�  b�$��HJ���џ �����+�=�O�a� s�����V���ͯ߯� ��'�9�K�]�o��� ��R���v�ؿ꿮�� #�5�G�Y�k�}Ϗϡ� �������Ϩ���1� C�U�g�yߋߝ߯��� ���ߤ��ȿ�<��� c�u��������� ����)�;���_�q� �������������� %7��@��d� P�����! 3EWi{�L�� ����////A/ S/e/w/�/HZl~ �/�??+?=?O?a? s?�?�?�?�?�?�?� OO'O9OKO]OoO�O �O�O�O�O�O�O�/�/ �/2_�/Y_k_}_�_�_ �_�_�_�_�_oo1o �?Uogoyo�o�o�o�o �o�o�o	-?�O _"_�F_���� ���)�;�M�_�q� ��Bo����ˏݏ�� �%�7�I�[�m���� P��t֟����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ 㿢��Ɵ(��O�a� sυϗϩϻ������� ��'�9���]�o߁� �ߥ߷���������� #�5���V��z�<�>� ������������1� C�U�g�y���J߯��� ������	-?Q cu�F�j��� ��);M_q ��������/ /%/7/I/[/m//�/ �/�/�/�/���? 0?�W?i?{?�?�?�? �?�?�?�?OO/O� SOeOwO�O�O�O�O�O �O�O__+_�/4?? X_�_D?�_�_�_�_�_ oo'o9oKo]ooo�o @O�o�o�o�o�o�o #5GYk}<_N_ `_r_��_���1� C�U�g�y��������� ӏ�o��	��-�?�Q� c�u���������ϟ� ���&��M�_�q� ��������˯ݯ�� �%��I�[�m���� ����ǿٿ����!� 3����x�:��ϱ� ����������/�A� S�e�w�6��߭߿��� ������+�=�O�a� s��DϦ�h������ ��'�9�K�]�o��� �������������� #5GYk}�� ���������� CUgy���� ���	//-/��Q/ c/u/�/�/�/�/�/�/ �/??)?�J?n? 02?�?�?�?�?�?O O%O7OIO[OmOO>/ �O�O�O�O�O�O_!_ 3_E_W_i_{_:?�_^? �_�_�O�_oo/oAo Soeowo�o�o�o�o�o �O�o+=Oa s������_�_ �_�$��_K�]�o��� ������ɏۏ���� #��oG�Y�k�}����� ��şן������ (��L�v�8������� ӯ���	��-�?�Q� c�u�4�������Ͽ� ���)�;�M�_�q� 0�B�T�f��ϊ���� �%�7�I�[�m�ߑ� �ߵ��߆������!� 3�E�W�i�{���� ����Ϧϸ����A� S�e�w����������� ������=Oa s������� '����
�l.� �������/ #/5/G/Y/k/*|/�/ �/�/�/�/�/??1? C?U?g?y?8�?\�? ��?�?	OO-O?OQO cOuO�O�O�O�O�O�? �O__)_;_M___q_ �_�_�_�_�_�?�_�? o�?7oIo[omoo�o �o�o�o�o�o�o! �OEWi{��� �������_>�  ob�$o&�������я �����+�=�O�a� s�2������͟ߟ� ��'�9�K�]�o�.� ��R���Ư������ #�5�G�Y�k�}����� ��ſ�������1� C�U�g�yϋϝϯ��� ��ʯ�����گ?�Q� c�u߇ߙ߽߫����� ����ֿ;�M�_�q� ������������ ������@�j�,ߑ� ������������! 3EWi(��� ����/A Se$�6�H�Z��~� ��//+/=/O/a/ s/�/�/�/�/z�/�/ ??'?9?K?]?o?�? �?�?�?�?���O�E�$FMR2_�GRP 1ZE�� ��C4  B�� 	� � VOhLS@Fw@ ~EE���B�~A�:{A�L�FZ�!D�`�D��� BT��@�{�ÖM?�  �O��<S@6����B���5�Zf5��ESQ�MA�  �_0[BHT�@JQ@_�33@�TPXSB�<RDx_�]S@@OQ��_�N�_�_RA<�z��<�ڔ=7��<�
;;�*߲<���M8����9k'V8���8���7�?�	8(���_?o �_<ouo`o�o�o�o�'�,B_CFG [9KThB�o/�i�NO 9J
�F0cq hp�lRM�_CHKTYP  )A� A@C@�0+A�ROM~p_MIN\�p�#���p�oP]X,@SSB�c\E TF���%�s���eTP�_DEF_OW � �$AC$�IR�COM�p5��$G�ENOVRD_D�O�v�!b�THR֥v d�dh�_E�NBT� h�RA�VC2C]�w�p �vE� ��o$��Lq2�C�fZ �ȁ�OU5@c9Lkq8fH9�fE<�p�O���d���ԟ��#C�  D+�1���L�\�@OAC�B�gAI�iI����ɀSMT2Cd�։E@�p'��$HO7STC�b1e9I�p���/R@ MC��$?����&�  27.0M�16�  e-�z��� ������h������:�ѿ˳	anonymous>�l�~π�Ϣϴ��"��Q@�� ��+�-��a�B�T�f� xߊ�Ϳ��������� ��K�,�>�P�b�t�� �����������5�� (�:�L��	������� ������� $6 H������������ ��� c�DV hz�������� �
//_q��� m/��/�/�/�/�/7 ?*?<?N?`?�/�� �?�?�?�?�?3/E/W/ i/k?\O�/�O�O�O�O �O?�O�O_"_4_WO �?N_|_�_�_�_�_O O+O�_?_0osOTofo xo�o�o�O�o�o�o�o o]_>Pbt� ��_�_�_��Go (�:�L�^��o������ ��ʏ�o�1�$�6��H�Z���ߡENT �1f��  P�!鏫�  �� ��֟ş������B� �N�)�w���_����� 䯧��˯,���b� %���I���m�ο���� �ǿ(��L��p�3� iϦϕ��ύ��ϱ�� �����G�l�/ߐ�S� ��w��ߛ��߿���2����V��z�=�QUICC0��c�u���1�����&���2�'���v�!ROUTERw�S�e���!PCJOG�����!192.�168.0.10����CAMPRT,��!1 >�%RT��BT� �!Softwa�re Opera�tor Pane�l�{�NAM�E !��!R�OBO0S_C�FG 1e�� ��Aut�o-starte�d�tFTP� ��ޏ����/ #/5/~�Y/k/}/�/� �/F/�/�/�/??1? �pw��|?�/��? �?�?�?�?�/O0OBO TOfO�?O�O�O�O�O �O�O����qOG_ �?�_�_�_�_�_�O�_ oo(o:o]_�_po�o �o�o�o�o__1_C_ Eo6y_Zl~�� eo�����1� D�V�h�z������o�o ���
�M.�@�R� d�v�9�������П� �����*�<�N�`�r� ��Ǐُ���ޯ!�� �&�8���\�n����� ��ǯI�ÿ����"� 4�w������������ ���������Ͽ0�B� T�f�xߛ�߮����� �����K�]�oρσ� t�Ϙ�������� ��(�:�L�o���������������_ERR g&�����PDUSIZ  �q�^���>~$WRD ?e�R��  guestq�dv�����SCD�_GROUP 3�he i{�I�FT$PAO�MP _�SHEDS $�CCOM��TT�P_AUTH 1�i <!i?Pendan���q�n1!KAREL:*����KC//'/��VISION SCET� �/\/m6!�/ �/�/��/�/�/�/7?�? ?m?D?V>�CT_RL j�8�q�
q�FFF�9E3y?P�FR�S:DEFAUL�T�<FANU�C Web Server�:�2R� L^�<YOkO}O�O�O��O��WR_CON�FIG k��?�?��ID�L_CPU_PC�@q�B�S�%P ;BHUMIN\�~)UGNR_IO���2q�	PNPT_�SIM_DO[V�e[STAL_SC�RN[V ��6oQT�PMODNTOL8�We[>ARTY|X%Q�jVy �ENB�W��
SOLNK 1l -o?oQoco�uo�o�obMAST�EZPijUOSL?AVE m�e�RAMCACHE��o�RO�O_CF1G�ocsUO� ~rCMT_OP@8]R
OsYCL�o+u��0_ASG 1n�G>
 �o�� ����*�<�N�`��r��������k�rNU�M1	
rIP��owRTRY_C�NZ+u�Q_UPD1,a� r8pr�o�n� g�� PR�CA_ACC 2�p�  W��� H��  ;�p 6� 6q�#�q���6��O������4̜�}�BUF001 �2q�= ���u0  u0�
���+�:�K��[�l�{�����u0�iH���u0�c`�� ���V������!��U0��A��P��a��Uq�����������U���Æ�҆�ㆤ������$��3�D�T�e��t��������u�������Z��������U'��6��G��V��Ug��v��������U������Ɇ�؆�	����2���$� )�-�)�5�)�=�)�E� )�M�)�U�)�]�)�e�<)�m�t� �t�)� }�~���������� ���¥��­��µ��� ����Š��͠��ՠ�� ݠ��堑������� ���������� ��%��-��5�� =��E��M��U�� ]��~�l��u��}� ҅�����ҕ��ҝ� �ҥ��ҭ��ҵ��ҽ� ��Ű��Ͱ��հ��ݰ���少�����s�#8�����3�� +�2�-�;�2�=�K�2� M�[�2�]�k�2�m�2� e���q񄣓Ú╢�� �⥢�Úⵢ�Ú�Ţ �Ú�բ�Ú���Ú� ��Ӛ�����#� �%�3��5�C��E� S��U�c���l�{� �}���\���Ӛ� �Ӛ򭲻Ӛ��Ӛ� Ͳ�Ӛ�ݲ�Ӛ���Ӱ�����q2r�� 4�<�5\\<�\PS]R}�HIuS�t� ܛ�� 2023-08-1�7+o��@���ΑR�\;��P5G|=Wk� �������� //0/gyf/x/�/ �/�/�/�/�/�/??/ Q/>?P?b?t?�?�?�? �?�?�??)?O(O:O LO^OpO�O�O�O�O�? OO __$_6_H_Z_ l_~_�_�_�O�O�_�_ �_o o2oDoVohozo h	�w���o�o�o +Sd%* d��Er0k�_�_ �o������� 1�C�U��������� ��ӏ���	��-�d� v�c�u���������ϟ ���<�N�;�M�_� q���������˯ݯ� &�8�%�7�I�[�m�� ������ǿ������ !�3�E�W�i�{ύϟ� h	��o�o�o���� ,�>�P�����RpC	 �ߗ�ѿ�������� �'�9�K�]�o�߸� �߷����������#� 5�G�~�������� ��������1h� z�gy����� ��	@R?Qc u������ */)/;/M/_/q/�/�/�/�/��I_CF�G 2u�� H�
Cycle �Time�Bu{sy�Idl2��min�+z��Up�&�R�ead7DoYw+8'? ;2�#�Count�	N'um �"����<���1�aPROG��"v����� �?�?O!O3OEOWO29��eSDT_ISO�LC  ��� ��@�.J23_D�SP_ENB  ��K80�@INC �w�M�Ø@A  � ?g�=���<�#�
�A�I:�o �A_(_��_P_��G�0GROUP �1x�KEr<A �C��_X_?��?�_��Q�_o!o�3o�_Woio{o�o��@_b[IN_AUT�O  ���J�@POSREC�C�b71��hKANJI_M�ASK�f�jKAR�ELMON y�˰?��yRok}�����.)r�3z�7��C���u�ouCL;_L�`NUM�@
���@KEYLOGG'ING�`����Q�E��0LANGUAG�E ��q���DEFAUL�T ���LG�!Y{�:72���x�@߰  880H [ ���'0�������cOy�;���
�(UT1:\�� ��.� @�W�d�v�����������(Z���LN_DISP |�O�48�_�_!�OCTOL`���Dz�0�A�A�v�GBOOK }��dޔz��ᑮ�Xٌү������,�<���83N�*�	 ��ۉ�QmK��aO�A���_BUFF 2~N�K ���235 ݿ������17�'�T� K�]ϊρϓ��Ϸ��� �������#�P�G�Y�����C��DCS ��9�B�AK�����%��� ��$��IO ;2��� !Z��Q�]�m���� �����������!�5� E�W�i�}����������������8�ER_ITM�Nd�ofx ������� ,>Pbt�����p�;SEVt�`�M7TYP�N�U6/H/Z/��aR�ST(���SCRN�_FL 2�F��0����/�/�/??(?:?k/TP>��O%"}M=NGNAM�D�ǥq���UPS)�G�I� 	��E�1_�LOADPROG� %g:%	T_ARCWELDG?��MAXUALR�M%��a� ��E
�B�1_PR�4�` h��L�@C,�����hO���%��ODoPP �2��� �ؖ	 %/�O�O�O�O_-__ Q_<_u_X_j_�_�_�_ �_�_o�_)ooMo0o Bo�ono�o�o�o�o�o �o%[F j������� �3��W�B�{���p� ����Տ��ʏ���/� �S�e�H���t����� ���Ο��+�=� � a�L���h�z�����߯ ʯ����9�$�]�H�DBGDEF �YE��eOu�_LDXDISA�0f;6�MEMO_AP�0�E ?g;
 ��F������/��A�S�e�@FRQ_�CFG �YG6��A F�@���H�<��d%h���yϋ���B�YKL��*�/� **:(�H��-���H� S�eߒ߉ߛ��߿��� ��J�YE'� �N�<�R�`�,(�ߥ��� ��������*��N� 5�r���k������������JISC 1�g9� �P�JL� ��`K���� �_MSTR ����SCD 1�ֽ��/�S>w b������� //=/(/M/s/^/�/ �/�/�/�/�/?�/ ? 9?$?]?H?�?l?�?�? �?�?�?�?�?#OOGO 2OkOVOhO�O�O�O�O �O�O_�O_C_._g_ R_�_v_�_�_�_�_�_ 	o�_-ooQo<ouo`o �o�o�o�o�o�o�ox;�MJPT��1��i�{�w^s�MIR 1���^�p ��Lx��.s< ���?O�.q?y�3\�N�� � ���P����.��©� &��5C��o.q ���~�+yH��@�b� ��v���Ə珺�� ��ҏD�b�4�^���b� ����П��؟�+y�� ��L�^�����g�q� ��ͯk�ů����� K�-�~�����5�W�ɿ ����׿ϯ��G�-� ?�a�c�q�����g�y� �������U�;�]� ��qߓ��ߣϵ��� �߽�?���3�=��a� ������������ J�\������e�w�� ��i���������I +�|��3U��� ���E+=�_�o^pKdq��j{  �\rLT�ARM_��ju�p�xtop/$^p�METPU  �.r���]qND�SP_ADCOLx3%�>.CMNTT/ G%FNp t/E'�FSTLI�/�'MST ���/xs�� ?
4G%POSC�F�'.PRPMls/9STR 1�j}=4�q<#�
�16q �5�?�7�?�?�?�?�? �?�?.OO"OdOFOXO �O|O�O�O�O�O_�A�G!SING_CH�K  �/$MOWDAQ��jy���@UDEV 	�jz	MC:t\HOSIZE3 ��@UTASK %jz�%$123456�789 �_�U>WT�RIfp�j{ lju%�8oh+oloOm��t�SYP�Q{uVT�?SEM_INF �1��XQ`)�AT&FV0E�0uo�m)�aE0�V1&A3&B1�&D2&S0&C�1S0=�m)A#TZ�o@'tHDl�a`o�#xA������ �oC��o ,��P���� ����֏?�Q�8�u� (�:���^�p������ ��)�`�M�����>� ����˯ݯ�����Ɵ ؟�[��������� h�ٿ�������3�� ��i��.�@�����v� ������пA���e� L߉ߛ�NϿ�rτϖ� �����=�O��s�&߀��R�������m_N�ITOR� G ?��[   	EOXEC1�"3�2:�3:�4:�5:�`<�U7:�8:�9:�5� �ҟ�9��E��Q�� ]��i��u����P������2��2��U2��2��2��2��U2��2��22�3��3��3E�@QR�_GRP_SV ;1��k (�A �o����MO�Q�_D��^�ION�_DBJP�N]�!�  �� �� ��gT?.@/L��20�20�gT��N� � �� �L�>cY-ud1�U�����aPL_NA_ME !e���!Defau�lt Perso�nality (�from FD)��aRR2� 1��L�XL�yx�hP d� W/i/{/�/�/�/�/�/ �/�/??/?A?S?e?@w?�?�?�?�?_X2F/ �?OO%O7OIO[OmOO�OaR<�?�O�O�O �O__'_9_K_]_o_��_���O�^
�_�_�P�_oo/o AoSoeowo�o�o�o�o �o�o�o�_�_O as������ ���'�9�K�]�, >������ɏۏ��� �#�5�G�Y�k�}�������� H�6� H�b H\���������d��"��E�S�Ő������������� ��ٯϯ��� �5�W���z������	`ï��Ͽ�>��:�oA!"���%�7� A�  Lɨ�'tw[k �����me~� �G��hȟ���ϰ����Ϡ���
�C��R� �1��u��@ � ����п @D�  ��?���Ӂ�?����A��6Ez  �Ѽ���;�	l��	� �@� 0v�w�� ���� �? � ��5��J��K ���J˷�J� ��J�4�JR�<�(�7'��d�5�@��S�@�;fA�6A��A?1UA��X@�O���=�N��f������T;f���X��5���*  ��  ß5��>������ҘM�?� ?�￰#������6�w�(� �>�5Ә��P�H��u�Uu�(y��u������5߫�N�	'� �� ��I� ?�  �Y�L��:�È��È=��������� <��� �� � ��e���?����@I�p�~�e���z��@!�p@�Wa�@��@��@��[C��C� �� ���B��C��d��@�7�  ���3�?���K�L͈����I�@�m�D �՚�������`(
%Y:a�� >�x?�ff0d�K/]/� ���/Ĥ+�8Y �/�*>���=��I���&���6)������_>��A!E�<2�!�<"7�<L���<`N<D��<��,-�j?y/������"I�?ff�f?m?&�0q�@�T싹1?�`�?Uȩ?X� �1W	�1������? ��O�7��|/QO<OuO `O�O�O�O�O�O�O�O_W�5FZ_S_ _w_�?�_Ij_�_fXHmN H[�YG� F���_ oo
oCo.ogoRo�o vo�o�o�o�o�et} �o`��_T�_{�o� ���t?���/� �S�>�w�b�U��Uɲ�Cq�֏m���������D�/�W	�ç��®�>�BH�� �� T��� ��x����@I�Y��@n�@���@: @l���?٧]�� ���%�n��߱���=�=�D��������@�oA�&{�C/� @�U����+J8��
�H��>��=3�H��_E� �F�6�G���E�A5F�Į�E��m�����fG��E���+E��EX�����>\�G��ZE�M�F�lD�
�п��� 
���.��R�=�v�a� ������п����߿� �<�'�L�r�]ϖρ� �ϥ����������8� #�\�G߀�kߤߏߴ� ��������"��F�1� j�U�g�������� ������B�-�f�Q� ��u����������� ��,P;t_� �������:%7p+�(-�4g�t-1���]3�ϩ�����4 �{������0+#���j�b/+/1E���|�0G+E)�/s/�/P�/�/�,.uPe2P�.q(?{4?^?I?�?m9F ��?�?�?�?�?�?�?��$OOLO 7OpO[O�O;?�O�O�O�Le�O�O1__A_g_U_1)m__�_�_�_�_�_j  2� H�6��H�,@",c\���B�������Bȓ���A��@ ��so��w��o�o�o�o�o-z#o5o,>TP`|���D������Aotc��
 `����� �&�8�J�\�n�����ؤ�#�rr���H�-��$MR_CABLE 2��(� V`2T*0aa@3 ?w��Lab��{�?`B?`�C �3!OM�`B����M�.�t �D�hr3&��J`�N`B�S`�O�
�v7��A�>�t D�UkA%W��i�Z`�J`CW`9�-��⋕�(ArrD��Z`���%*!��S` �C�/��7 7�����<|�cD����� �Z�+u�M�_�į�� ͯ�����ݯ�T�O� %�q�I�[����ɿ7��!���(�:�1(�pi�{ύ�1(*���** ݃OM }����HV s�W�%% 2345678901�ς�� ����3  � jba3 3!
����not segnt ��?�W�%�TESTFE�CSALGRPgD0*bad�ԈqF�
��0�0k~h������1(9UD1�:\mainte�nances.xsml�_�  �z��DEFAU�LT�l݂GRP {2���  p�t�g3%  �%1�st mecha�nical chgeck�3!���#����U� �j�7�I�[�m��3"��c�ontrolleAr��������T(����!3E��MX��m3""8�3 ���U������P
C��3�W�������ڔ�C��ge��. battery�G/�U	tI/[/m/�/�/��Supp�ly greasXQ�/����#<��!�/�U8/??1?�C?U?���cab!l�/�/�?,(
�/�? �?�?OO�����?�?��?�O�O�O�O�O%@$�O_Ը׿4_ �OY_k_}_�_�_�O �__&_8_�_o1oCo Uogo�_�o�_�_�_�o �o�o	jo�oQ�o @�o�����0 ��f;��_�q��� �����ˏ�,��P� %�7�I�[�m������� �ǟ�����!�3� ��W�������ܟ��ï կ���H��l�~�S� ��w����������� 2�D��h�=�O�a�s� ��Կ����
����� �'�9�Kߚ�o߾��� �Ϸ���������N߶� 5��$��}���� �������J��n�C� U�g�y��������� ��4�	-?Q�� u���������� f;��q� �����,/P b7/�[/m//�/�/ ��//(/�/L/!?3? E?W?i?�/�?�/�/ ? �?�?�?OO/O~?SO �?�?�?�O�O�O�O�O 2O�O_hO_�Oa_s_ �_�_�_�O�_�_._o R_'o9oKo]ooo�_�o �_�_�oo�o�o#85�l�b	 TCp ���o����� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=��  ��a?� ; @�a �x� �����fd�ɯۯ�hw*�** �a �f��?�A�S�e�'���8���������o�c $�¿�"�4���X�j� |�ƿؿ�P������� D��0�B�Tߞϰ�� �߮���
ߔ����� d�v߈�&�t���Z��������*�<�j�$�MR_HIST �2��e;�� 
� \�b$ 2345678901K�(S���J�9�o�� ��s����o(�� ��^p�9K�� �� �$6�Z ~�G�k�� �/�2/D/�h//��/�/U/�/ �SKCFMAP  �eW>���z �z �/�%ONREL  z$;��!�� �"EXCFEN�B%7
�#�%>1FN�CE?74JOGOVLIM%7d;�0�"WKEY%7�5�5_PAN$8�2�2�"�RUN�<�;SF?SPDTYPe805��#SIGN%?74TO1MOT�?41�"�_CE_GRP 1��e�#C�[p ���Oz#|O�O&D�O�O �O__�O>_�ON_t_ +_�_O_�_�_�_�_o �_(o�_Lo^oEo�o9o �o�o�o�o�o�o�o�6�k�!QZ_ED�IT"D�'CTCO�M_CFG 1���-H5��� 
�vq_ARC_B2�%Ep9T_MN_M�ODE"F�P9U?AP_CPL�T4�NOCHECK {?�+ �/ S�e�w��������� я�����+�=�O��a�;NO_WAI�T_L!GkwV@NTF~q��+�ez#��o_ERR`A2��)�!���
��.���1PS�e����pOᓫ��| H��+q�K��p��@D�����`£�9��!\�x)<�0�� ?�k�Яk��0��ڒPARAM:⒬�+�O�,�S�>��!p��� =  ����������ۿ�ɿ ��#�5��Y�k�G�=���ϯ�B���BODRDSP�s$FP8�OFFSET_C�ARap$�	�DIS���S_A�pAR�K"GlyOPEN_FILE5�$A�qlv��pOPTION_�IO�?�1��M_P�RG %�*%$�*����i�WOU�-�fGP���	�z$��   2P�#�9��#�	 �x(#���z#���RG_DSBL  3���!̚����RIE�NTTO$0z!Cٴ0�!A ��UT�_SIM_D����"P���V��LCT ���hr�q�zz%d��_PEX ��8�+�RAT � d�P5+��UP )���|��������Rz ��z z Y2�1���$�2_C��L�XL�x��%��� +=Oas��� ����'9 K]o�z'2� ����
//./@/ R/ã�|/�/�/�/�/ �/�/�/??0?B?�il&k/|>��|?�?ϒP�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�?�?_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo�O�OTofo xo�o�o�o�o�o�o�o ,>Pb��Co�=����}!��� ��~����}�}��W�B�{�.�$�p��� ������ҏ؏���n�`��<�K�I�p�	`���~�������:�o�����ҟ�����A��  �i�'��.j����a��me?b �������e���q�������@�˯�������Os��1����� ��l�@ �]��G� @D7�  Z�?�`�F��?��b���D�  �Ez|�Y5�  ;��	lr�	 ��@�� 0g�h��� ��V�� � �� �в��H0�#H��G��9G�ģG�	{Gkf���S�X�,���C��\��%�D	� D@� D��	�������  �5��>�t�[�ù�b�tφ� �B��Bp{����!����O�^�#�8��� а���������6���U:�(:��:��]��T���p��	'� �� ��I� ?�  ���=��Ͳ���^�߶� <���� � � �*�^��u�"^��5���N��\�&���t�?���C��C	����B[���J��x��i0Z��@������������������
�@��2�v���_� \�G���k��������Ә������:!��>�x?�ff%�"�� [�Wi���8���
>�� �n���IкX�����������$�>����
�<2�!<"�7�<L��<`�N<D��<���,�/>`����
�?fff?�2�?&l��@T���~?�`?U?ȩ?Xǎ�9 ��gs���b��`�� P��A//:/%/^/ I/�/m/�/�/�/�/�/ �/?�/6?���/?��?+8HmN H[����G� F���?�?�?�?O�?,O OPO;OtO_OqO�O�E 9��M�O%�S?_w?@_ �Od_v_�_�_9�_�_�[_�_�_oo<o'o ���fb�wkC6o�ox2o�o�m?���o��o	�o��çs��Tsm��H�����Z�d��`�a�q@I�܊�@n�@���@: @l��?٧]j� ��%�n��߱���?=�=D�ɺ�p���@�oA��&{C/� @��U� �+�J8��
H���>��=3H���_
� F�6��G��E�A�5F�ĮE���2�D���fG���E��+E�?�EX�Z�D��>\�G�ZE��M�F�lD�
[���iϏ��� ޏ��;�&�_�J�\� ��������ݟȟ�� �7�"�[�F��j��� ��ǯ��į���!�� E�0�i�T�y�����ÿ ���ҿ���/��,� e�Pω�tϭϘ��ϼ� �����+��O�:�s� ^ߗ߂ߔ��߸����� � �9�$�I�o�Z�� ~��������������5��r(�q4��9����j�"�3��ϩZ�l��q4 ��{�����q�0+#8������jb����1E�䴛|[ 
	J8n\��J�EP*P��A�O �@��#G2 �MT�x����r$��/�5/ /�Y/ �O�/z/�/�,e �/�/�/�/?,??�A)2?D?z?h?�?�?��?�:  2 H��6�vH��3\Ŵ�vBoacao`B�XpWpA�p@so8OJO@\OnO�O�O�M�CP/@�O�O�O__%\�v�N$�p�p�A84T�3�u
 %__ �_�_�_�_�_�_�_o�!o3oEoWoio�z7R�����H-��$�PARAM_ME�NU ?
��  �MNUTOOL�NUM[1�w��`F�`�`�iA�WEPCR�`.$�INCH_RAT�E�`SHELL�_CFG.$JO�B_BASp �WVWPR.$�CENTER_R�Ir�`$tAZIM�UTH OPTB��a$tELEVATION TC�a�$tDWqTYP�E SNqARCLINK_AT(p?STATUS�c�y�__VALUq��`LEP�a.$WP_�`�b��|�� ���$�6�_�Z�l��~����aSSREL?_ID  �����USE_PR_OG %�j%��<���CCRTƄ���c�_HOST !�j! �]��AT� '�y�@�R�{�����_TIMEO�U$��g  �`GDEBUGƀ�k���GINP_FLM3SKޟ�TR��[PG�p  ���O�L�CH��yr�k�@����ү����� �C�>�P�b������� ��ӿο����(� :�c�^�pςϫϦϸ� ������ ��;�6�H��Z߃��WORD �?	�k
 	sRS;�ZPN�q�[MAIp��S�UNq��TE��Z�STYL5r��CO�LX�
��L� U �U�0�d��TRACECTL� 1�
�a� � Q ��I�D/T Q�
��d�D � ������������7P�� UP��p���MP��IP�⨿���������	���
��U�������������0�B�T�������ȀZ�l� ��� �����������@@@�@@@@*@@@0	 &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO`�O�O�O�MI�LEp�ȁ]P�`�=�I�_�UP ��[P8Y��q ���NQY��}d�bG_zj��zj��&�_DEF�SPD ��k2�Ђ  Т`I�NPTRL �����a8dU�QPE__CONFIP�X��̈́}aw $�L�IDS��� 	gL_LB 1�X�m���dTB�  B4Vc}fn�Obljio�e�W_ << ρ?��k�o�o�o�o  �o6NlR�d�����ZZ o��=�4�a��fQ�C�𠏓�ď
eGRP �1�;l�,�@�  �[�_aA�?x�D P�D?V�C2���k��E�d-�=��Qw �}���o&aY�´��r�[�B�����������П����_a>'oY>a���K�]��G� =N�=R�b���^���ѯ�� ���z��=� �M�s�^�  Dz����_`
��ɿx�ٿ���#� �G�2�k�VϏ�zό�@�ϰ������j�)Q�
V7.10b�eta1_dN �B(�A�\)�A�G���F�>��^���F�Aw���n�ffF��A�p�AgaG��q�q@�����V� ߳�������_cAp@�
�U`�#� 5�G�BҢQ����� z��v�����F�B�ga���Ru0��e:� �@+�a��QG�@���l�� B{PB���z�BH������� ���g��;Q)��
�x��xR�N�0n��P��R{ �w���W�qd�KNOW_M  ��e+VdSV �����U ��I[m��|�P�_b5�
cMރ��`�V�	BU����3/�CTߞ��?��@ {Q{�{Pr%n/�,�pa+MRރ��T�כּ�
��/�+̍OADB�ANFWD�+cS�Tށ1 1�Y84�Uk�V�l?_V T?f?x?�?�?�?�?�? �?�?;OO,OqOPObO �O�O�O�O�O�O_�O__572@<	!S?_`G�<}_Q_߀3g_y_�_�_574�_�_�_�_575oo1oCo57A6`oro�o�o577�o�o�o�o578*�<57MA 06��ds�WOVLD  �\{,/ȏ72PARNUM  C;���63SCH�y �u
B��P�.3b�UPD��um����U_CMP_��p���/',5ĄER_wCHK҅��,10"�Ϗ�RS� #?N�_MO ?C�_0�~�U_RES_G?0�\{
��]����� ֟���+��0�a�T� ��x���������fP����Я���P��� ��`,�K�P���_`k� �������`��ɿο�� p��υ�Xp(�G�<Lυ�V 1�F�P�	!@[l�F�T?HR_INR� �q��,5d��MASS6�� Z��MN�����MON_QUEUE �\u,6S��U�TNɀU�N
�3�J�ENDO�m�i��EXEx�iՎ�BE�w�Y�J�OPTIO�V�v�M�PROGR�AM %-�%�LІ�1�K�TASK�_I�t��OCFG� �-��!�T�D�ATA��]�~��2%�������� ���/�A�S�e�w�"������������INFO�ǡ�<ԍ�* <N`r���� ���&8J@\n������ȡ�c ��S�I�K_W���]��ENB��p�[Q&2/(G�W�2�� X,�		�=���&j/�%�!$N0���)�)���_EDIT �]��/�/P�WERFL�خ�23�RGADJ �^�*A�  55?���A5��6M���\u��?�  Bz3W��<�!����%n�?8�/W3�2Y�c7�	HD�l�ǩ��p1?� Ax�ɻt$F*%@/'B **:0B��#O�5CQM\ujBeE��AoI���?�O]M �MmOO�O�O�O/_�O �O__!_�_E_W_�_ {_�_o�_�_�_�_�_ soo/o]oSoeo�o�o �o�o�o�oK�o5 +=�as��� #��������9� K�y�o���������� ۏ�g��#�Q�G�Y� ӟ}�������ş?�� ��)��1���U�g��� �������ӯ���	� ��-�?�m�c�u�￙� ��ٿϿῦ�	p�z� �0hϡό�I��C����ϋ��&�S7PREOF �c:�0�0�
5IORITY����&�1MPDSaP��:���UT?�|C6ODUCT<���*)��6OG�_TG0A��*���HIBIT_DO�	8�TOENT �1��+ (!?AF_INE��^�~�7!tcpi�>��!ud���?!icm��>���XY\3��,��1)� =A�/��0��X�;�G���k� ������������&@8\C��*��\3�c9��?���3�>w�7�=G/�GL�9�4��8�>A~�2,  �YЀ�����5�6)Z)�
//./�3��ENHANCOE ճ�2A�Ad(�/u%��B��J��\�11PORT�_NUM���0�x�1_CART�REP���S2SK�STA��+�SLGmS[�����3��0Unothing�/s?�?�?�<Y?��?�?�?��61TEM�P ����?8���0_a_seiban��bO��rO�O�O �O�O�O�O_�O(__ %_^_I_�_m_�_�_�_ �_�_ o�_$ooHo3o loWo�o{o�o�o�o�o �o�o2BhS �w������ �.��R�=�v�a��� ����Џ���ߏ���<�'�`�O61VER�SI������ �disable��"KSAVE ����	2670/H755J�]����!~/�����/� 	�S���:�I�|��e@��¯ԯ���J����.�9����_�� 1���|�T��������;�URGEbM B �$���WFİ ��h"��WW�崖���*WRUP_DE?LAY �>ص�R_HOT %�_Ƹ�}/e���R_NORMALD���T�<��x�SEMI�Ϯ�|��9�QSKIPd�	ܺ'u�x[�2�W�V� h�z�=�Gš߯י��� ���߹���'�M�_� q�7��������� ����7�I�[�!�� m��������������� !3EU{i����G��$RBT�IF�
<RCVT�MOU75��� DCRd���� �I�A�3��B��B3��@��5@�7��*�=������~�����T �rL���N=ߍ�� �<2�!<"7��<L��<`N�<D��<��,��V���-  /)/;/M/_/q/�/�/��/�/�/�/�/��RD�IO_TYPE � k���/EDP�ROT_CFG ���2��BHfͳEE9
�2�W;7 ��B�j0�? �:��?��?�?OM �?KO��rO�ߓO��O �O�O�O�O_�O5_CW aOf_�-_�_}_�_�_ �_�_�_�_�_1oS_Xo w_yoo�o�o�o�o�o �o�o=oBaou ������� �9>�]��_��� ������ݏˏ�#�(� :���[����m����� ��ٟǟ���$�C�� W�E�{�i�����ï���ӯ	�/� ��G7INOT 2�Gɔ1�AG;� ^�p��2�<��
Hf�0 ��Ȼ ��ٯ�����B�0� f�L�vϜϊ��Ϯ��� ������>�,�b�t� Zߘ߆߼ߪ������� ��:�(�^�p�V�� ����������� ��6��EFPOS1� 1�9  x�)c3������ ��*�w�����$H ��l�+��a ���2D�� +�w�K�o� ��./�R/�v// �/�/G/Y/�/�/�/? �/<?�/`?�/]?�?1? �?U?�?y?OO�?�? �?\OGO�OO�O?O�O cO�O�O�O"_�OF_�O j_|__)_c_�_�_�_ �_o�_0o�_-ofoo �o%o�oIo�o�oo�o �o,P�ot� 3��i���� :�L���3������ S�܏w� �����6�я Z���~������O�a� ����� ���D�ߟh� �e���9�¯]�毁� 
����ɯ�d�O��� #���G�пk�Ϳϡ� *�ſN��rτ��1� k��Ϸ��ϋ�߯�8����5�n��Z�2 1�f��"�\������� �"��F���C�|�� ��;���_������ ��B�-�f����%��� I��������,�� P����I��� i���L� p�/�Sew �/�6/�Z/�~/ /{/�/O/�/s/�/�/  ?�/�/�/?z?e?�? 9?�?]?�?�?�?O�? @O�?dO�?�O#O5OGO �O�O�O_�O*_�ON_ �OK_�__�_C_�_g_ �_�_�_�_�_Jo5ono 	o�o-o�oQo�o�o�o �o4�oX�o Q���q��� ��T��x����7� ��[�m������>� ُb�����!�����W� ��{����(�ß՟� !���m���A�ʯe�� ���$���H��l��x��v߈�3 1�� =�O�����+�1�O� �s��pϩ�D���h� �ό�߰������o� Zߓ�.߷�R���v��� ��5���Y���}�� *�<�v��������� ��C���@�y����8� ��\�����������? *c���"�F� �|�)�M� �F���f� �/�/I/�m// �/,/�/P/b/t/�/? �/3?�/W?�/{??x? �?L?�?p?�?�?O�? �?�?OwObO�O6O�O ZO�O~O�O_�O=_�O a_�O�_ _2_D_~_�_ �_o�_'o�_Ko�_Ho �oo�o@o�odo�o�o �o�o�oG2k� *�N����� 1��U����N��� ��ӏn��������� Q��u����4�������4 1���j�|� ��4��X�^�|���� ;���֯q�������� B�ݯ��;������� [���ϣ��>�ٿ b�����!Ϫ�E�W�i� �����(���L���p� �mߦ�A���e��߉� �߿����l�W�� +��O���s������ 2���V���z��'�9� s�����������@ ��=v�5�Y �}���<'` ���C��y /�&/�J/��	/ C/�/�/�/c/�/�/? �/?F?�/j??�?)? �?M?_?q?�?O�?0O �?TO�?xOOuO�OIO �OmO�O�O_�O�O�O _t___�_3_�_W_�_ {_�_o�_:o�_^o�_ �oo/oAo{o�o�o  �o$�oH�oE~��=�a�П�5 1�ퟗ��a� L������D�͏h�ʏ ���'�K��o�
� �.�h�ɟ��퟈�� ��5�П2�k����*� ��N�ׯr�����Я1� �U��y����8��� ӿn�����϶�?�ڿ ���8ϙτϽ�X��� |�ߠ��;���_��� ��ߧ�B�T�fߠ�� ��%���I���m��j� ��>���b������� �����i�T���(��� L���p�����/�� S��w$6p� ����=�: s�2�V�z ���9/$/]/��/ /�/@/�/�/v/�/�/ #?�/G?�/�/?@?�? �?�?`?�?�?O�?
O CO�?gOO�O&O�OJO \OnO�O	_�O-_�OQ_ �Ou__r_�_F_�_j_��_�_o��6 1���_�_o�oyo�o �_�oqo�o�o�o0�o T�ox�7I[ �����>��b� �_���3���W���{� �����Ï��^�I��� ���A�ʟe�ǟ ��� $���H��l���+� e�Ư��ꯅ����2� ͯ/�h����'���K� Կo�����Ϳ.��R� �v�Ϛ�5ϗ���k� �Ϗ�߳�<������� 5ߖ߁ߺ�U���y�� ����8���\��߀�� ��?�Q�c������"� ��F���j��g���;� ��_����������� fQ�%�I� m��,�P� t!3m��� �/�:/�7/p// �///�/S/�/w/�/�/ �/6?!?Z?�/~??�? =?�?�?s?�?�? O�?xDO*o<d7 1�Go �?O=O�O�O�O�?_ �O'_�O$_]_�O�__ �_@_�_d_v_�_�_#o oGo�_koo�o*o�o �o`o�o�o�o1�o �o�o*�v�J� n���-��Q�� u����4�F�X���� ޏ���;�֏_���\� ��0���T�ݟx���� ������[�F����� >�ǯb�į����!��� E��i���(�b�ÿ ��翂�Ϧ�/�ʿ,� e� ω�$ϭ�H���l� ~ϐ���+��O���s� ߗ�2ߔ���h��ߌ� ��9�������2�� ~��R���v������ 5���Y���}����<� N�`���������C ��gd�8�\ ��	���c N�"�F�j� /�)/�M/�q/WOiD8 1�tO/0/ j/�/�/?/0?�/T? �/Q?�?%?�?I?�?m? �?�?�?�?�?PO;OtO O�O3O�OWO�O�O�O _�O:_�O^_�O__ W_�_�_�_w_ o�_$o �_!oZo�_~oo�o=o �oaoso�o�o D �oh�'��] ��
��.���� '���s���G�Џk�� ���*�ŏN��r�� ��1�C�U����۟� ��8�ӟ\���Y���-� ��Q�گu��������� ��X�C�|����;�Ŀ _�������Ϲ�B�ݿ f���%�_��ϫ��� �ߣ�,���)�b��� ��!ߪ�E���i�{ߍ� ��(��L���p��� /����e������� 6�������/���{��� O���s�������2���V��z��/�$M�ASK 1�+����XNO�  ���MO�TE  �$G_?CFG �N���PL_RAN�GJ?�%��OW_ER �%���SM_DRYP�RG %�)�%�K��TART ��	*UME_�PRO��e/�$_�EXEC_ENB�  ?�GScPD> � �(�(gTDB�/�*RM�/��(IA_OPTI�ON����!_AIRPUR�� F*B?�M�T_� T�L��`1g�o=�"C�?  N?�?�?�?��??1OBOT__ISOLC�>0�~zENAME� F*T/�	OB_CATEG�� �O�DuCO�RD_NUM ?��;1H?755  ?�O��OY� PC_TI�MEOUT� x�� S232g1���# LT�EACH PEN�DAN!Pc�pT��=JH Mai�ntenance_ Cons?m_�?"�_DNo Use�=�__�_�_�oo%o�9RNPO� #R�56QC7H_LA �?� �	�aso!UD�1:�ouoR� VA3IL�A5�1_SR  /;1���eR_INT7VAL6��Yp�> yV_DATA_GRP 2��� D>pP �����y�!� �A�/�e�S���w��� �����я���+�� O�=�_���s�����͟ ���ߟ���K�9� o�]���������ǯ� ۯ���5�#�Y�G�i� k�}�����׿ſ��� ��/�U�C�y�gϝ� ���ϯ��������	� ?�-�c�Q߇�uߗ߽�������$SAF�_DO_PULS�K�A? ��CSCA�NR6�<@SC����`�X�!? �1
�2��A�Q�U
[�? ����� ������|��#�5�G�XY�k�Hrc�2��[��d����>9	X�Hi @��� ��?��. �p�_ @3�T01n���YT D����� ��"4FXj |������Bo�Le���Vp,/>/F$
*  iU�;�o�Tg!Eqp�duE
�t���Di�@�k�Z  � �+Jk���A S��/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_�_�_.a����_�_�_ oo)o;oMo_o�_�� �o�o�o�o�o�o�o	 -2qoo0�"�# �%�-~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N��_r������� ��̯ޯ���o8� J�\�n���������ȿ 3auk���,�>� P�b�tφϘϪϼ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{�@��������(�� ����/�A�S�e�w� ��������������+=��
�T�.�����"z��	123456�78�"h!B�!���������f��'9 K]o��	��� ���//(/:/L/ ^/p/�/�/�/�/�/�- ��/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO�/�/TOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_3O�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �_�o $6HZ l~������ �� ��oD�V�h�z� ������ԏ���
� �.�@�R�d�v�5��� ����П�����*� <�N�`�r��������� ̯�����&�8�J� \�n���������ȿڿ ����"����DςV��{ύϟϻ
�Cz  Bp�� �  ���2��� } 6���
���  	���2<�#�5�G�Y�i���j��߯��� ������	��-�?�Q� c�u��������� �����)�;�M�_�q� �������������� %7I[m�B�� j�k����<�� ��  ������
�>
�t  ��
�"��`�$SCR�_GRP 1��*P30� �� ��� ���	 m�u� k����ǒ���ί�����C� ��݌*'����LR Mat�e 200iD �567890��LRMc# 	L�R2D j ��
O1234i%�x�,m�� �&_u��@d�d�ӻ����)	�"?%?7?I?�[?k<��H�u�$yd�?��? �?�?�#����?(O�?LO�>K� h���,W��  [d�B���ƗOȕB�D�A���O  1@���E�@��@�O# ? �E�BH��_��J�F@ F�`8R@_7Od_O_�_s_ �_�_�_�_�_o��A��AR1oo.o@oRdB�`o�_�o�o�o�o�o �o�o$H3lW �~ߥz#��w���A�������A@ O>��,��@�@4U����k��'�,�;ϫ���A�@�v΅$�?�5ۀ���"��A ��*��z�M�HY�k�:�h���
�� ����ß��ҟ����Y/k#DECLV�L  ������"܂A��*SY�STEM*��V9.10214 s��8/21/202o0 A � `��o�SERVEN�T_T   $� $S_NAM�E !��PO�RT����ROT�O�� ��_SPD���J�B�̠T�RQ   
^ɣAXISҡק�Ϡ 2 �ɣDE�TAIL_ � l $DAT�ETI����ERR�_COD(�IMP�_VEL�� 	�:�TOQB�ANGwLESB�DIS���N���G��%$LI�N(���ɣREC�ҡ ,�����F�MRA�� 2w d��IDX��܊�ߠ h�$�OVER_LIM�I���	��OCC�URҡ  �-�COUNTER��� �SFZN�_CFGҡ 4� $ENABL�(�ST"���FLA�G��DEBUF�R[� ���Jҡ� � 
$MI�N_OVRD���$I��W�{�s���F�ACE�|�SAF>��MIXED�̄��d�{�ROB��$�NE��PPôHE�LL �	 w5$J��BAS(��RSR_.�  ?$NUM_�B�� �1w��2�9�39�49�59�6�9�79�8w�	�RO�O��~�CO��ON�LY�p$USE�_AB���AC�KENBA���IN�۰T_CHK��O?P_SEL_9���g_PU���M_%�;OU��PNSֽ����x�9���M3�TPFWD_KAR@���.�RE��$O�PTIONX�$QSUE 鿠D;�Y���$CSTOPI_3AL����EX����l��(�XT��M1���2��MA��STY���SO��NB��DI��TRIFÄ�@�INI��Mà��NsRQ���END���$KEYSWI�TCH'�<����H}E=�BEATMo�PERM_LE?�RG�E<�n�U;�F���<�S��DO_HO�M��O����EFP0����G��STL���C��OM)���OV�_MS�ѻ�ET_IOCMN�Ӕ����]���HK��
 gD -Ǳ�SU'�f��MP��.�PO�¿$FORC&�W�ARNOM� ��@$FUN�C� 7�U���ART���2�3�4~T]��OL�Lo���!�UNLO�%���ED%��p�S�NPX_AS#�; 0$�ADDV�X��$SIZ(�$�VARw�MULTKIP���� Ao � $�� ��	&�� ��'�yC;�kFRIF���۰Sl�~	��[NF��ODBUS_A�D�&ү���CM�1�DIA]$D�UMMY1���3��4��SО�� � X�TEt���8�SGL#!�TA��  &�8�<#'�� 5 $ ST�MT��U#PSEG̵�U!BW��%$SHsOW]%��BANi OTPOF��9�i0���ȠVC���Gh� 1 $PCp�ܰ� �$FBk-P�(SP��A���%��VD� g�7� � �A0��0� b�$1� +7� +7� +7T� +75)96)97)9U8)99)9A)9B)9@} +7�+7r +7F)8 � �859��8O9	 �8�i91v91�91�91��91�91�91�91
�91�91�9���G59U2B92O92\92i9U2v92�92�92�9U2�92�92�92�9U2�92�93(9359U3B93O93\93i9U3v93�93�93�9U3�93�93�93�9U3�93�94(9459U4B94O94\94i9U4v94�94�94�9U4�94�94�94�9U4�94�95(9559U5B95O95\95i9U5v95�95�95�9U5�95�95�95�9U5�95�96(9659U6B96O96\96i9U6v96�96�96�9U6�96�96�96�9U6�96�97(9759U7B97O97\97i9U7v97c�7�97�9U7�97�97�97�9e7�97�4��VPk�=UТ ٠���.�
����� x? $TORu��+  D�M��RΠ��ߔQ_��R��P��G B�S��C=��F'�_U� 2�Z��a��Lu��� �  �3ǚ
J�$0��<^��"VALU3����A�����FO�ID_YL���HI��I]?$FILE_�����$��M�SA�ϱ hҐ�E_BLCKo�#�>!>,�D_CPU<� <�
>����J�x���R  � �PW���В��LA�c!Sα������R?UN_FLGŵ�� ɱ��?�̵걡�걬��Hิ���]�T2�A�_LIo � �G_O���I�P_EDI�� 1$���,�4��	���7�]�#�BC24 � ��̰� ��,�FT�����TDC̰A��C���aM�������TH�"S�����R��� . ERVE�������������� �X -$:�L�EN��G���:в�R1Ak��N�W_�i�i1:�פ2��MO4��S���I��#��0��Ք:о�DE�ա�LACE���CC8�#��_MA� ��8����TCV�/���T!�0�O�E�2��P�!s����!J��A�%�M�䟠J�0������F�2���� ������ JK��VK@�!��������J�!l���JJ�JJ�AAL��1��1�+�d
!/�5��b�N1V�Pb�!��!�L��_Q!؞�1��CF� =`ҐGROU��?!���!N��CS��R�EQUIR�E�BUj6љ�$T��2��7������ Ά� \w f�AP�PR��CL!�
$:=�N0CLOr�@	�S��U	�՜�> �n�M���a���'_MG�� C0�p�0	�BRK�	�NOLD�� RTCMO+��
��J+��P3���������PO���X���6 7 �1!7 �� ��a��!���PATH�����f؟� ��%�� S�CAj��1�INF9�UC�Д��C0KUM(Y������ 	!á�$*�$*:$ �PAYLOA�J{2L��R_AN��e#L��o)k!_){!��R_F2LSHR	Ԩ!LOp$��'#|�'#ACRL_y� �� �W$Y�H��!��$H�2FLE�X3 ��J�� P�ϧ�� �
�|409�  :F� X��Щ7�4[�Z���d�v߈�F1�1E"G��@�߻�������RBE�� ��1�C�U�g�y�� )XFT�����6@XX����1��T�W'QX �����D}H���U�H ����0�4�=�+�O�`X�j�|���R�BJ��! �����������Ƭ�AT;F���ELP�@{�s��J�� ��;JE� CTR�6A�TNƑ	v��HAN/D_VB!�31��nt" $�PF2�����SW�������~#� $$M � �	���x��|�@�u�vAƠ\ �šD��A����
A�AA���U��
D��D�P�G����S�T����	��N�DY˰. ��t�} ;� �'�1�'�!^'��}T�0�P�P(1:CL�U^g4�J��$ �p�4� �p��b���ASYM�#�����#���!�_ ��(�$����x/-/?/Q/c#Jj,|*p�����)HD_VIds�٨b�V_UN K�ؠ�� c�!J��� E���,��%(�L��-����)�/?���Sd$4,4 20��HRt��i�%zrͱF0@�D	I� ��O�}�ΰ�c�& 0`�I�A �#�<@'�'�?@|��20�@ϰ ' �[ �qME�At`hB�)�T�PT� �`�j����E0a��oȊ�~�T���� �$DUMMY1�:$PS_9@RYF�0ư$��� 7FLA��YP�S���r�$GLB_T`�p���j�N1T�wA:qF�( X ��t�ST�A��SBR��M21_V��T�$SV_ER� O���@�X�CL�@�A��@O�ɰGL�E�W��) 4��t�+$YqbZqbW������!�sAC�"�b��U.��* �PN�Ѕ��$GIJp}$�� )n�ѼЎ��+ L����S�}�$FS�E��NEA�R�@N@CF-�@T�ANC@B 
 JO�G�0 ,��?$JOINT�Q�P{ ��MSET��-  ��E�A�`�S�bȱ���`��.�� BpU�A?����LOCK_FOx� �q�BGLV=s�GL��TEST_sXM3 ��EMPi��PR�����$U�0���P2*���!�+��p��!�)B�C�E����B� $KA�R�AM�TPDRqA��_�V�VEC�0�p�Z�IU!�,&�H=E��TOOLC���VDREw�IS3�5��6C6@ACH|���-��O�rôĵ30a��SI# � @$RAIL__BOXE�Qe�oROBO��?�e�?HOWWAR1<����ROLM��7��a��H�a��*@vO�_F�`!e�HT'ML5��hr��t��w/b��Rz��O�20��0k�o �����OU~�1 d���))�r�a���$PIP��N �P������H@!� �0?CORDED���L� *�XT� ��)ɰ��`O)� 2 D ��OBE�s���P?����?S�qS;YS?ADRqɰ�j�TCH�p 3� ,�PENҲO1A���_����a'�
���VWVAE�4� � e����P�REV_RTR��$EDIT�VSHWR�a,� �BJ��٠DT��1'$~ a$HEADd�h��A t��KE�Ѿ��CPSPDX&JKMP\L�20R�@F�5GD1�I��5SrC^pNE��q�TwTICKC�M�M1ڐ�%HN"�6� @I�!�e`!_GqP�&��P0STY���LO��҂"�"��07 t 
�G��%$���=,�S`!$��PY�������P��&SQU�Y��5��ءTERC�n��ј�S�d8 ��8��g�P�g%Q��b�`Oo�b�D@IZ��4������PR%���B�!� PU�aE_�DO2�XSz�KN�AXI<@[&�UR�`�Cr � jd�q�`_��|ET}BQP��Xҕ;0Fҗ�<0A߁Ց��9���)��=�SRqt9l�0�y�R�z�E �v
Y�r�E�w�C��C �>U3�>UC�>US�PU@j]��PU�\��nYC�_�|]C�]L�^�p���� �0SC�� : he�DS� `��3SP�jeATA��r�A� �"��ADD�RES��B�SH�IF�c�_2CH�pfIмa�TuU�I�q ;��CUSTO�D8V
��I�<���~aC*��
��
�V�-ANG�= \*���;0|�1�0IrC��2�B�z�^�Iq�TXS�CREEA>ٰW1TINA{��Мt���}!~A~b��? T�![�B|Z�7��v�JA{JB�t�RRO��G�{R �q8���UE�$@ �ꐕ��9S|�|RSM� @G�U.�0�S�ͰS_ ��s��c�v����~A�C��O��t 2?�pUE��A�kҶ��@GMT_�L9��YAG�Ol��BB�L_��W��G�B ��;0�O���L�E�b*� �b)�RI;GH3�BRDmԤaOCKGR��[�T/|Z�W�WIDTH�� aB������2�I&j EY~`F�C�z �6 2��	ABAC�K1��Εq�M�F�O�LAB(Q?�(M�I����$UAR��0��S�H	�� D 8��G�_@!�b1�T�R�����C����B�O�aG�E�� x�T�U?��R��BLUM�aF�`GERV�S৐P1�j��FK��@GE�0�@5I LPѥ�B	E�0/a)�?a��Oa�������5��6��7��8ޢ�2b�@1�]tԳ�����S�0EUSR��G �<*�S�U���c��F�O�`��PRI�Amx��m�аTRIP��m�UNDO�H��`0�BE)AE����{@u0 I�,���AG H0T0[ a�a'�OSr�<�AR�@�Û�ӁJ��@�ӫ�c��$ˁ�U١ӁKl�~ό�٢�%çOFF����L(���O��"�Je����-Ke�GUvP�m�p�a)׻�SUB�"LtТ�RTe��DM�"�F�g �3OR��o�RAU�@p�T�٢U�9_��$N |�@��OWN��$S#RC���^0D�����BMPFI4a}@ESPA�2�p�����.!���� ��
 ӁO� `��WO$P���1�0COP��$r@�_�м�i��p�WA�C��M�#�L�1���5�a �P�rSHADO�W^@���_UNS�CA~�㓔��DGyD��WEGACc�w�VC P)�ӁQ� ��@l3$�ER�p,��1�����C� ,�DRI5V�6�A_V� O��� 6 D|�MY_UBY{�4�B6c�l5���0�p.!��1���P�_��4��L#KBMv&�$� DEY�cEX �'�t�MUv 1X&�h�US]�h@˰_R�q�����`����G�PPACIN�!i0RG��Xn��`n��n��i�REF���ac���n�RS �`[�Gt�PrH� ��RS��S���x����O�	h�:ARmE+SWf _Ag�� @O���aA(�`'�BEl�U.0H���[��HK32Tu�?���A$�pp�EA� zL�3�'A�C�MRCVӁU� �ʠO?0M3�Cs	��ð�REF��������C � ���!�!�1%�f_��|g(�xPSi����1�ˀ�ЄV �2�����04�����0OU�'�<�&4� Q�a�2��$�p_p@���S}ca�!D��`UL6�pT(�COG�H�3U 0NT#�P4�1�O5`�[6��[30L���5��5`��7����VIA_L�]`W� ��@HD�`Ɛ�$JOg����?$Z_UPL̰ �ZEPW�5�139����_LIM�$EP 1I�4��1�1�q�a���`Q%�6�X� �0}c�A@` }cCACH*LO!lD�A� �I��|���C@M%I�cFA�ETVP�FN�+$HO3���p@OCOMMJ�O�O=� �G�'��d3��͡�$ ��VP�p�6R_SI	Z*@TZR ;X�1<W��n�MP`ZFAIj�0Gl�@AD�Y�i�MRE�$�REWG�PU� ��s�ASY�NBUFs�VRTaD�U�TEQn�OL�`�D_��
eW��PC&�`TU �@QD�U�ECCU�VEM�� �ERb�GVIRC��Qe�SN��Q_DE�LA����簶�AuG�YRXYZ��}�W��h!�d��2o`T�IM�af��b���EGRABBJ`�Y+ PEЄY.�ڒLAS���PA_GEWEZ>���sbc_uT�#���)���I�t��fb�BG2/�V��p�PKq �f,XA�'GIOpN�)A�	��@�Q:�[����AS�P}FN�� LEXPv\��ӳ��z�Q��I �S��E���E���m��a��
��]��+��DY���\��*�ORDıȠ�p°@��"�^ $0TIT�ɰ�������VSFv���_�  ��$�[1 URl��1SM�`�����ADJ΀�0Z�D�a D��AA�L�0�PΠ
BPER�I<@��MSG_Qc$FQdU5���eBa�b���0�@���@��W�XS�h�c���� K�CH)�H�OL�� ���XVR�d7r+�T�_OVR2��ZABC\�e�6��C��
�0c�z�VS�@ f � �$_��|�CTIVz��AIO���FY��IT
�mDV	��
mX@��{Q��&àPS�!�� �S��p�A� ���ALSTY���A�00��_S���� Z�DCS;CH��g Lg�#��w��@ �GÀ@� EPG�NA�C���A"�_GFUN��@GqZ&�2�h���$L���}�qZMPCF\Ցi���
�����LN �.�
����`]�?j $�Az^��CMCM` Cr��C\����P^� O$J��D+Q !�2�+ǚ07Ś0Ǩ���0�c�UX�a��UXE&���a&�z�<��z����Ɍ����FT�F<1!����ٰ�Gk D�����
���Y@Dp l �8cR�PU��$�HEIGHY�?(0ؖ�����$�m � �S�$�B0A���L�SHIYFvS��RV@F�����+�C�0�\�-4��D��ְ^s�� UD,���CE��V}!Y����PHERh� �n ,00�F�X��r���FA;1��c����۠�S�HOT�_���@S�MIPOW�ERFL �pc�zk� ��WFDO`�� ��G@� 1 ������� L{!��_EIP����c��j!AF�z0E_�$���!F�T��S��w�!��x����f���!�R'`MA@�����@�����p��������[!OPCUA�\�
J�!CTPz0p���d���!
PM��X	Y��e�?��	�f.�!RD%M�V��gz��!R90�	�h�#/!
���@X�yi/o/!RL�P�Cp/�)8^/�/!�ROS���,�4��/?!
CE� M�T�@?�k�/S?!E	2C{�q?�lB?��?!2WASR�C��m�?�?!N2USB�?�n�?>7O!STM��QO�o&O�O���O�tO��M��I
�KL ?�%�� (%S?VCPRG1�OZ"U2__P3@_E_"P4h_m_P5�_�_"P6�_�_P7�_�_"P8ooP90o5kT�]oQ
_�oQ 2_�oQZ_�oQ�_�o Q�_%Q�_MQ�_ uQ"o�QJo�/Q so�/Q�o�/Q�o=� /Q�oe�/Q��/Q; ��/Qcݏ/Q��/Q �-�/Q�U�WQ��O �BG`�O P���'Q� ���1��U�@�y�d� ������ӯ������ �?�*�Q�u�`����� �����̿���;� &�_�Jσ�nϧϒϹ� �������%��I�4� m��jߣߎ��߲��� �����!�E�0�i��J_DEV ��?�MC:t��?GRP 2��b���@bx 	�/ 
 ,��q��� �������9� �2�o� V���z����������� #
G.k}�� �X����� 1U<y`r� ����	/�-/� "/c//�/n/�/�/�/ �/�/??�/;?"?_? q?X?�?|?�?�?�?�? F/O%OOIO0OmOTO fO�O�O�O�O�O�O�O !__E_W_>_{_b_�_ �_O�_�_�_o�_/o oSoeoLo�opo�o�o �o�o�o�o+=$ a�_V�N��� ����9�K�2�o� V�������ɏ���ԏ �#�zG�Y�@�}�d� ������ן������ 1��U�<�y���r��� ��ӯ�<�	���-�?� &�c�J����������� �ȿڿ���;�"�_� q�Xϕ�쯊��ς��� ���%��I�0�m�� fߣߊ������������!���W��d �^�	E��y���������	�%�	�.������G���G�W� e�O���s��������� � C���-Q? acu����� �)M;]� ������/� %//I/�p/�9/�/ 5/�/�/�/�/�/!?c/ H?�/?{?i?�?�?�? �?�?�?;? O_?�?SO AOwOeO�O�O�O�OO �O7O�O+__O_=_s_ a_�_�O�_�_�_�_�_ �_'ooKo9ooo�_�o �__o�o�o�o�o�o# G�on�o7�� ������aF� ��y�g��������� я'�M��]���Q�?� u�c����������#� �����'�M�;�q�_� ��ן�������ݯ� �#�I�7�m�����ӯ ]�ǿ���ٿ���� Eχ�lϫ�5ϟύ��� �������M�2�D��� ���eߛ߉߿߭��� %�
�I���=�+�M�O� a��������!�� ��9�'�I�K�]��� ������������ 5#E�������k �����1s X�!���� ��	/K0/o�c/ Q/�/u/�/�/�/�/#/ ?G/�/;?)?_?M?�? q?�?�?�/�??�?O O7O%O[OIOO�?�O �OoO�OkO�O_�O3_ !_W_�O~_�OG_�_�_ �_�_�_o�_/oq_Vo �_o�owo�o�o�o�o �oIo.mo�oaO �s���5� E�9�'�]�K���o� ���̏�������� 5�#�Y�G�}������ m�ןş����1�� U���|���E�����ӯ ������-�o�T��� ���u�����Ͽ��� 5��,���߿Mσ� qϧϕ������1ϻ� %��5�7�I��mߣ� ����	ߓ�����!�� 1�3�E�{�ߢ���k� ����������-��� ��z���S��������� ����[�@�	s ������3 W�K9o] ����/�#/ /G/5/k/Y/{/�/� �//�/�/�/??C? 1?g?�/�?�?W?y?S? �?�?�?O	O?O�?fO �?/O�O�O�O�O�O�O �O_YO>_}O_q___ �_�_�_�_�_�_1_o U_�_Io7omo[o�oo �o�_o�o-o�o! E3iW��o��o }�y���A�/� e�����U������ я���=��d��� -���������ߟ͟� �W�<�{��o�]��� ������ۯ���˯ �ǯ5�k�Y���}��� ��ڿ�������� 1�g�Uϋ�Ϳ���{� ����	�����-�c� �ϊ���S߽߫����� ����kߑ�b��;� ����������C� (�g���[���k���� ������� ?���3 !WEg�{��� ���/S Ac����y� �/�+//O/�v/ �/?/a/;/�/�/�/? �/'?i/N?�/?�?o? �?�?�?�?�?�?A?&O e?�?YOGO}OkO�O�O �O�OO�O=O�O1__ U_C_y_g_�_�O_�_ _�_	o�_-ooQo?o uo�_�o�_eo�oao�o �o)M�ot�o =������� %�gL����m��� ��Ǐ��׏��?�$�c� �W�E�{�i�����ß ������՟���S� A�w�e���ݟ¯��� ������O�=�s� ����ٯc�Ϳ���߿ ���Kύ�rϱ�;� �ϓ��Ϸ�������S� y�J߉�#�}�kߡߏ� �߳���+��O���C� ��S�y�g������ ��'���	�?�-�O� u�c������������ ��;)Kq�� ���a���� 7y^p'I# �����/Q6/ u�i/W/y/{/�/�/ �/�/)/?M/�/A?/? e?S?u?w?�?�??�? %?�?OO=O+OaOOO qO�?�?�O�?�O�O�O __9_'_]_�O�_�O M_�_I_�_�_�_o�_ 5ow_\o�_%o�o}o�o �o�o�o�oOo4so �ogU�y��� �'�K�?�-�c� Q���u����ҏ䏛� �����;�)�_�M��� ŏ���s�ݟ˟�� �7�%�[�������K� ����ٯǯ����3� u�Z���#���{����� տÿ�;�a�2�q�� e�Sω�wϭϛ���� ��7���+߽�;�a�O� ��sߩ�����ߙ�� ��'��7�]�K���� ����q���������#� �3�Y������I��� ����������a�F X1y������9]g�$�SERV_MAI�L  g]�~COUTPUTR_h @G�RV 2�  ` (�-�G�SAVEsaTO�P10 2� d c/+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_���YP�DFZ�N_CFG �`$��~MQGRP 2WW�� ,B   �A�PgD;� B}�P�  B4#�RB21�H7ELLPR	��Ħ�nW ok%RSRoo"o[oFo ojo�o�o�o�o�o�o �o!E0i{�~?�  �]r�����r� h ���r�q�x�r2h d��|�}8��VHK 1
�[ �r�|� v���ɏď֏��� �0�Y�T�f�x�����������\OMM ��_��RFTOV_ENBR��P��OW_REG_U�I0�EIMIOFWDL�����Ue�/WAIT-�1�oRȍ�mQ����TI�MQ���įVA�Q��e�_UNIT�,����LCJ�TR�YQ��GMO�N_ALIAS k?e���he �������úm���� 
��ǿ@�R�d�vψ� 3ϬϾ������ϟ�� *�<�N�`�߄ߖߨ� ��e�������&��� J�\�n���=���� �������"�4�F�X� j����������o��� ��0��Tfx ��G���� �,>Pbs� ���y�//(/ :/�^/p/�/�/�/Q/ �/�/�/ ??�/6?H? Z?l??�?�?�?�?�? �?�?O O2ODO�?hO zO�O�O�O[O�O�O�O 
_�O_@_R_d_v_!_ �_�_�_�_�_�_oo *o<oNo�_ro�o�o�o �oeo�o�o�o8 J\n�+��� ����"�4�F�X� �|�������]�Ï� ����ɏB�T�f�x� ��5�����ҟ����� �,�>�P�b������ ����g�����(��ӯL�^�p�����>���$SMON_DE�FPROG &������� &*SYS�TEM*��߷�p��?��REC�ALL ?}��� ( �}9co�py frs:o�rderfil.�dat virt�:\tmpbac�k\=>169.�254.E�120:4504߿d�v����}0�mdb:'*.*/�A� K������ ߓ�4x�:\ ��$е�����`�r߄� }5�a"�4��� P�������*ϳ��� _�q���1��L��� ���ߧ߹�J�[�m� ���#�5��������� �"��F�Wi{�� ��;������� ��B�Sew����- ��R��,� �a/s/�/�3/�N/ �/�/?��/L]? o?�?�%?7?��?�? �?/$/�/H/YOkO}O �/�/=O�/�O�O�O?  ?�?D?U_g_y_�?�?�/_�?�_�_�_�Lx�yzrate 124 �_�_�_[omo�o�D!h:n170�8�@=oOo�o�o }:O,O�o�bTfx�K1�O5�kL� ���[�_5o�g�a��s���}6�_+�=� �Q��􏇏tpdisc 0���b���ˏ\�n����Ctpconn 0 ;� 5�G�؟���!� EV�h�z���:�� ԯ�������A�ӯ d�v�����,�>�Q��4����
f1 ���� ɿZ�l�~ϑo�o�oG� �������!���E�V� h�zߍ���:�ï���� ����0�A���d�v� ����,�>�Q������ �+ߴ���`�r����߀2���M��������$SNPX_AS�G 2����%� � 0�%�M � ?�PARAoM %/� �	;P�r�P��& � OFT_KB_?CFG  �+�OPIN_SI�M  %���( RVN�ORDY_DO � ��:QS�TP_DSB���~SR �%	 � & �LAB_WELD3_1�����TOP_ON_E�RRG�PTN� % ��A	"RING_�PRM�YVCN?T_GP 2��2 x 	zy/�`g/�/�/�/VDN �RP 1u	�  �!%�/�/?#?5?G? n?k?}?�?�?�?�?�? �?�?O4O1OCOUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�_�_�_oo )o;oMo_o�o�o�o�o �o�o�o�o%L I[m���� ����!�3�E�W� i�{�������؏Տ� ����/�A�S�e�w� ��������џ���� �+�=�d�a�s����� ����ͯ߯��*�'� 9�K�]�o��������� ɿ�����#�5�G� Y�k�}Ϗ϶ϳ����� ������1�C�U�|߀yߋߝ߯������"P�RG_COUNT���"��ENB�4/��M$��1�_U�PD 1�T  
���{��� �����������/� X�S�e�w��������� ������0+=O xs������ 'PK]o �������� (/#/5/G/p/k/}/�/ �/�/�/�/ ?�/?? H?C?U?g?�?�?�?�? �?�?�?�? OO-O?O hOcOuO�O�O�O�O�O �O�O__@_;_M___ �_�_�_�_�_�_�_�_�oo%o��_INF�O 1i�9O�q`	 Ho�o�wo�o�i?���@Cz=��oޝk���?a³?����33�o�`��� A�e @� p>�@ >����k C��7���$���6��B �p4?q��vL��KzrC3����Sp B�3����YSDEBU)G	�j��?`dR�zpSP_PASS	��B?�{LOG �ffs�  2?`�hEo  �aq`�  UD1:�\�tLn�r_MPC �}i�:�L�i��bk��i��SAV ��y�a�q�r;e� �SV�TEM_TIME 1�wt� 0?`����;cʇMEMBOK  i�N��p��N�`�p�X|�O�� @p�;c�@����ǜ�������q �k@�0�B� T�f��o��������ү�;c���!�3�E�@W�i�{�������e�� ӿ���	��-�?�Q� c�uχϙϫϽ�����`����)�̅SK%��*��9�i�{ߍ߁��:?`4,�2�����A��p��?a ֒" ��� ��$�T�f�x�<l���� ����Ԁ��������	����݀�+�P�b�t�����?`$ ����������, >Pbt���� ���(:.��T1SVGUNS�PD�u '�u��]2MODE_LIM ,����}�f��}XAS�K_OPTION�p-���_DI~�pENB  ����u�BC2_GRP 2LՌs�%/�֑�C�9#QBC?CFG +��c ���/t&`�/ �/�/�/�/�/ ?? D?/?h?S?�?w?�?�? �?�?�?
O�?.OO>O dOOO�OsO�O�O�O�O�O_;d�L _�OS_ e_�OB_�_�_�_�_�_ q�o/��Po1ooUo Coyogo�o�o�o�o�o �o�o	?-cQ s������� ���)�_�E�0Ps� ������ǏE��ُ�� !��E�W�i�7���{� ����՟ß����/� �S�A�w�e������� ѯ�������=�+� M�O�a�������q�ӿ ���'ϥ�K�9�[� ��oϥϷ��ϗ����� ���5�#�E�G�Yߏ� }߳ߡ���������� 1��U�C�y�g��� ����������ѿ3� E�c�u���������� ����)��M; q_������ �7%[Ik ������� //!/W/E/{/1��/ �/�/�/�/e/?�/? A?/?e?w?�?W?�?�? �?�?�?�?OOOOO =OsOaO�O�O�O�O�O �O�O__9_'_]_K_ m_o_�_�_�_�_�/�_ o#o5oGo�_koYo{o �o�o�o�o�o�o�o 1UCegy� ������	�+� Q�?�u�c��������� ͏Ϗ���;��_S� e�������%�˟��۟ ��%�7�I��m�[� �������ůǯٯ� ��3�!�W�E�{�i��� ����տÿ����� -�/�A�w�eϛ�Q��� ������߅�+��;��a�O߅�o֣��$T�BCSG_GRP� 2o���  �� 
? ?�  ���� �����(��$�^�H�Ђ��Ү���d�@ ���?��	 HBL������?B$  C�����	�����Cz	�Q�A�Д�333?&f�f?����A�����a� ���͘��|���DH����@��q��t� ����D"w�����d/
 ��r����u������:I�c	V3.00~��	lr2dI	*�}�ҔS3 � ���  �/+��J2����fG/$%�CFG !o�e�� ��K*�u"q�x,�,��/ �/�*x��/�/�/?	? B?-?f?Q?�?u?�?�? �?�?�?O�?,OO<O bOMO�OqO�O�O�O�O �O�O�O(__L_7_p_ �_�����_�_�_[_�_ �_�_oo>o)oboMo �o�o�o�owo�o�o �o:�я�_k�o q������� %��5�[�I��m��� ��Ǐ��׏ُ�!�� E�3�i�W���{���ß ���՟����5�G� �g���w�����ѯ�� ����+�=�O��_� a�s�����Ϳ߿�� ��'��K�9�[�]�o� �ϓ��Ϸ�������� !�G�5�k�Yߏ�}߳� �����������1�� U�C�y�g���Y��� ������	�+�-�?� u�c������������� ��;)Kq� �O����� 7%GI[� ������/3/ !/W/E/{/i/�/�/�/ �/�/�/�/??A?S? ��k?}?;?9?�?�?�? �?O�?OO+OaOsO �OCO�O�O�O�O�O_ _'_9_�O]_K_�_o_ �_�_�_�_�_�_�_#o o3o5oGo}oko�o�o �o�o�o�o�oC 1gU�y��� �_?��!��Q�?� a���u�����Ϗ��� ��)��M�;�q�_� ������˟������ %��I�7�m�[�}��� ��ǯ���ٯ���� !�3�i�W���{����� տÿ����/��S� A�wω�3��ϳ�9�o� ������=�+�M�s� aߗߩ߻�yߋ����� ��9�K�]�o�)�� ������������ 5�#�Y�G�i���}��� ���������� UCyg���� �������EW /u����� /�)/;/M/_//�/ q/�/�/�/�/�/?? �/7?%?[?I??m?�? �?�?�?�?�?�?!OO EO3OUO{OiO�O�O�O �O�O�O�O�O_A_/_ e_S_�_w_�_�_i�_ �_�_�_+ooOo=o_o aoso�o�o�o�o�o��o'K9oY~ s �p�s �v���r�$TBJO�P_GRP 2"�au� / ?��v	�r�s�$�|�ip��@� �0�u  � �� � � �=�t @�p�r	 �BL  I�?Cр D�w�q�e�>�n�j�|�<��B$?����@���?�33C�S���a���ǇI�[�x}����;�2�������@��?���z;���V�A�g��〝 ���6�ƕp>̧�����;���pA:�?�ff�@&ff?�ff��ޟa� ��u�󄦁x��,�:v,���c?L����ʐDH�x^�d�v�@�33�����>ʐ������8���퉡�q=�2�D"�����������x=�9�K�9��ݯ ﯐�������חɿ�� ��� �����?�Y�C� Q�ϰϋ�E�������0���@ߙsC��v2����	V3.0~�	lr2d�t�*���t�q�ߤ�� E8� EJ�� E\� En�@ E�pE�� �E�� E�� �E�� E�h �E�H E�0 �E� Eϻ���� E��� �E�x E�X �F���D�  �D�` E���P E��$��0���;��G��R��^op Ek��u�����І��(��� �E��Н�УX O9�IR]�)�q��������v���9�՟���tESTPARSr��x�p�s�HR��ABLE �1%�ys��tD��� `��������w�q��	��
�����.��q�������t��RDI��q-�?�Q�c�u�����O��	%7HI[�S���s �� .@Rdv�� �����//*/ </N/`/r/�}� ��r ,��)����~�������������"NUoM  au�q%��p s�t��_CFG &�;�/3=�@�pIMEBF_TT��*5�s���6VERr��!�6��3R 1'� �8�ߙr�p7A dp�/  O1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_�_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[���� �����!�3���RA_|1�6@�5��MI_CHAN�7� �5 ��DBGL�Vڀ�5�5�ᡀE�THERAD ?U������G��E����血ROUmT�0!�
!S��q�D�SNMASK���3��255.���wӭ���џw���O�OLOFS_DI���k�ӉORQC?TRL (Kg��O�T>�s������� ��ͯ߯���'�9� K�]�o�������=�ƿ������PE_DE�TAIǈ�PGL�_CONFIG �.�9�1��/�cell/$CID$/grp1�@d�vψϚϬ�b�:� ��������1���U� g�yߋߝ߯�>����� ��	��-����c�u� �����L������ �)�;���_�q����� ����H�Z���%7I�.}��������G1ۿ�� ��6HZl~��� �����/�2/ D/V/h/z/�/�/-/�/ �/�/�/
??�/@?R? d?v?�?�?)?�?�?�? �?OO*O�?NO`OrO �O�O�O7O�O�O�O_ _&_�OJ_\_n_�_�_ �_�_E_�_�_�_o"o 4o�_Xojo|o�o�o�o Ao�o�o�o0B�=��User� View R�}�}1234567890s����`��t^�2����Yy2fy�o7�I�[�m������`r3�ߏ���'�9���Z��4 Ώ������ɟ۟�L���5��G�Y�k�}� ���� �¯�66��� ��1�C�U���v��7꯯���ӿ���	�h�*��8��c�uχ���ϫϽ������ �lCameradzZ�#�5�G�Y�k�}�[Eߧ߹��� q����	��-�?�5�  ���ߏ��� ���������1�|�U�g�y���������� ��͉F���1C U��y������ ��	������� gy����h� �	/T-/?/Q/c/u/ �/.��[� /�/�/�/ ??/?�S?e?w?�/ �?�?�?�?�?�?�/�� 驊??OQOcOuO�O�O @?�O�O�O,O__)_ ;_M___O�����O�_ �_�_�_�_o�O)o;o Mo�_qo�o�o�o�o�o r_��Q�bo);M _qo��������%�7��o�g9 �x���������ҏy ����+�P�b�t�P������9�	��00� ���	��-�?��c� u���.�����ϯ�� ������۩�^�p� ��������_�ܿ� � K�$�6�H�Z�l�~�%� ��r�������� �� $�˿H�Z�l߷ϐߢ� �������ߑ�˕���� 6�H�Z�l�~��7ߴ� ����#���� �2�D� V����J������� �������� 2D�� hz����i�� �+Y 2DVh ������� 
//./��"K�z/ �/�/�/�/�/{�/
? ?g/@?R?d?v?�?�?A-  E)�?�? �?�?O#O5OGOYOkO<}O�K   �?�? �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� ��������L�  
A (  }�0( 	 � G�5�k�Y���}����� Ïŏ׏���1��U�:��J ��/�� ����1?�����*� <�C#��f�x���џ�� ��ү����O�,�>� P���t���������ο ����]�:�L�^� pςϔ�ۿ������� 5��$�6�H�Z�l߳� �ߢߴ����������  �2�y�V�h�z��ߞ� ����������?�Q�.� @�R���v��������� �����_�<N `r������� %&8J\� �������� /"/4/{X/j/|/� �/�/�/�/�/�/A/? 0?B?�/f?x?�?�?�? �???�?OOa?>O PObOtO�O�O�?�O�O �O'O__(_:_L_^_ �O�_�_�_�O�_�_�_� oo$ok_K�@  FbSoeowoFcMg1����+frh:\�tpgl\rob�ots\lrm2�00id�`_ma�te_�b.xml 3o�o�o%7I0[moV���� ������,�>� P�b�t��������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l��� }�����Ưد����  �2�D�V�h��y��� ��¿Կ���
��.� @�R�d�{�uϚϬϾ� ��������*�<�N� `�w�qߖߨߺ����� ����&�8�J�\�n�:�h�Q Mo�`�<< �` ?�n��n�������� �/��G�e�K�]�� ���������������3aoV�$T�PGL_OUTP�UT 1yQyQ/ ���� ����0B Tfx����� ��//,/>/P/�����f 2345678901u/�/�/ �/�/�/�#oRr/�/? "?4?F?X?�/\?�?�?�?�?�?n:}�?OO ,O>OPO�?�?�O�O�O �O�O�OxO�O_(_:_ L_^_�Ol_�_�_�_�_ �_t_�_o$o6oHoZo loozo�o�o�o�o�o �o�o 2DVh  ������� �.�@�R�d�v���� ����Џ�􏌏��*� <�N�`�r�������� ̟ޟ�����8�J� \�n����q}�ᶯ@ȯگ����!�@���E�W��� ( 	 Z/��z�����Կ ¿����
��R�@� v�dϚψϾϬ����� ����<�*�`�N�p�@r߄ߺߨ���h&��� �����*��L�^�8� ���b*������q��� �����C�U���Y��� %�w���������	g� ��?��+u�a� ����); Gq����S ����%/7/�[/ m//Y/�/}/�/�/�/ I/�/!?�/?W?i?C? �?�?�/�?�?�?�?O O�?%OSO�?;O�O�O 5O�O�O�O�O_eOwO =_O_�O[_�___q_�_ �_+_�_o�_�_9oKo %ooo�o�_io�oQo�o �o�o�o#5�ok }�����G Y�1��9�g�A�S� �����ӏ��я�����Q�c���)WGL1.XML!�����$TPOFF_LIM ��+�������N_�SV��  (����P_MON M2��+�+��2��STRTCHOK 3���������VTCOMPA�T՘_�ĖVWVA/R 4����ٔ� 6� ��������_DEFP�ROG %$��%
LAB_WE�LD_1����_D?ISPLAY��$��ʢINST_MSwK  � �?INUSERU���LCK^�%�QUI�CKMEN���S7CRE����`�?tpsc�^�м�����Ұ_ֹST�S���RACE_C_FG 5����u��	��
?��?HNL 26٪��A��� ��uχϙϫ������������IT�EM 27a� ��%$12345�67890H�Z� � =<R�xߊߒ� G !�ߠ۬�\� �ߣ�F��j�*�<�� R����ߟ��ߺ���� ��v�f�x����(� ��~��������>�P� b�����2Xj��v ����L �*�����  ��6�Z�5/� P/�`/�/�/��/ / 2/D/�/h/?:?L?�/ p?�/�/�/|?�?.?�?  Od?O�?�?cO�?~O �?�O�OO�O<ONO_ rO2_�OB_h_�O�O�O __&_�_J_�_o.o �_Ro�_�_�_To�_�o �o�oFo�ojo|o�o `�o���o�0 �T�x8�J��`� �$����ȏ,�؏�� �t��������6��� ����ğ(��L�^�p� �����f�x�ܟ�� � �ۯ6���Z��,����B���Ư���S'�8|-ϔ��  �Ɣ� 9���
 �����B�úUoD1:\O������R_GRP 19�5�� 	 @렚Ϭ˖��Ϻ������ޠ$�;�I���O�s�^ߗ߂�?�  ���ۮ�������� ,��<�>�P��t����������(�	�b�<�N���SCBw 2:�� �� �������������*��UTORIAL ;��6�u���V_CONFIG <��4��2����OUTPUT �=��� �� �$6HZl~� ������� $/6/H/Z/l/~/�/�/ �/�/�/�/�// ?2? D?V?h?z?�?�?�?�? �?�?�?	?O.O@ORO dOvO�O�O�O�O�O�O �O_O*_<_N_`_r_ �_�_�_�_�_�_�_o _&o8oJo\ono�o�o �o�o�o�o�o�oo" 4FXj|��� �����0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� ��P�b�t����� ����ο����(� �L�^�pςϔϦϸ� ������ ��$�5�H� Z�l�~ߐߢߴ����� ����� �2�C�V�h� z������������ 
��.�?�R�d�v��� ������������ *;�N`r��� ����&8 I\n����� ���/"/4/EX/ j/|/�/�/�/�/�/�/ �/??0?A/T?f?x? �?�?�?�?�?�?�?O O,O>OO?bOtO�O�O �O�O�O�O�O__(_|:_����Y_ k_UQD_�_9��_�_�_ �_oo&o8oJo\ono �o�oEO�o�o�o�o�o "4FXj|� ��o������ 0�B�T�f�x������ ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߽߬� ��������*�<�N� `�r��������� ����&�8�J�\�n�����������$TX�_SCREEN �1>mUUP�}�����	-?Q���V��� �����bt! 3EWi{�� ����//�A/ �e/w/�/�/�/�/6/ H/�/??+?=?O?�/ s?�/�?�?�?�?�?�? h?O�?9OKO]OoO�O �O
OO�O�O�O�O_ #_�OG_�Ok_}_�_�_�_�_<_�_�$UA�LRM_MSG k?����� �_ ��o-o^oQo�ouo�o �o�o�o�o �o$�H�USEV  �
mzv�RECFoG @�����  ��@�  }A�q   Bȶ�
 I������ ��%�7�I�[�m��������qGRP 2�A�{ 0��	 ����PI_BB�L_NOTE �B�zT��#l������p���DEFPRO`%
k (%<c��� Q���u�����ҟ���� ��,��P�;�t���FKEYDATA� 1C��Ӏp 	�w��֏ٯ�¯�!���,(-�T����(POINT � ]\�^�WEL�D_ST������P���߿��END N���TOUCHU�P��  ORE INFO8�;�x� ��qϮϕ�������� ��,�>�%�b�I߆ߘ�� ��/fr�h/gui/wh�itehome.png�������������point��S�e�w���*����arc_strA�E�������'�{���weldB�]�o�������4���enK�����(��touchup��@ew�������wrgA��� /��8\n��� �E���/"/4/ �X/j/|/�/�/�/A/ �/�/�/??0?B?�/ f?x?�?�?�?�?O?�? �?OO,O>O�?POtO �O�O�O�O�O���O�O _ _2_D_V_]Oz_�_ �_�_�_�_c_�_
oo .o@oRo�_do�o�o�o �o�o�oqo*< N`�o����� �m��&�8�J�\� n��������ȏڏ� {��"�4�F�X�j��� |�����ğ֟����� �0�B�T�f�x���� ����ү������,� >�P�b�t���������ο��ϟ��}������:�@L�^�6πϒ�l�,~� ��v��������A� (�e�w�^ߛ߂߿��� �������+��O�6� s�Z��������� ��O'�9�K�]�o��� �������������� ��5GYk}� ������1 CUgy��,� ���	//�?/Q/ c/u/�/�/(/�/�/�/ �/??)?�/M?_?q? �?�?�?6?�?�?�?O O%O�?IO[OmOO�O �O�ODO�O�O�O_!_ 3_�OW_i_{_�_�_�_ @_�_�_�_oo/oAo �eowo�o�o�o�o�_ �o�o+=O�o s�����\� ��'�9�K��o��� ������ɏۏj���� #�5�G�Y��}����� ��şןf�����1� C�U�g����������� ӯ�t�	��-�?�Q� c�򯇿������Ͽ� 󿂿�)�;�M�_�q�  ϕϧϹ�������~� �%�7�I�[�m��V`����V`����߼��ݦ������,��3���W�>�{� ��t���������� ��/�A�(�e�L����� ����������  =$asRo��� ��� �'9K ]o����� ���#/5/G/Y/k/ }//�/�/�/�/�/�/ ?�/1?C?U?g?y?�? ?�?�?�?�?�?	O�? -O?OQOcOuO�O�O(O �O�O�O�O__�O;_ M___q_�_�_$_�_�_ �_�_oo%o�_Io[o moo�o�o2o�o�o�o �o!�oEWi{ �������� �/�6S�e�w����� ����N������+� =�̏a�s��������� J�ߟ���'�9�K� ڟo���������ɯX� ����#�5�G�֯k� }�������ſ׿f��� ��1�C�U��yϋ� �ϯ�����b���	�� -�?�Q�c��χߙ߫� ������p���)�;� M�_��߃������h�����p����p����,�>��`�r�L�,^��V ����������!E W>{b���� ���/S: w�p����� //+/=/O/a/p�/ �/�/�/�/�/�/�/? '?9?K?]?o?�/�?�? �?�?�?�?|?O#O5O GOYOkO}OO�O�O�O �O�O�O�O_1_C_U_ g_y__�_�_�_�_�_ �_	o�_-o?oQocouo �oo�o�o�o�o�o �o);M_q�� $������� 7�I�[�m���� ��� Ǐُ����!��E� W�i�{�������ß՟ �����/���S�e� w�������<�ѯ��� ��+���O�a�s��� ������J�߿��� '�9�ȿ]�oρϓϥ� ��F��������#�5� G���k�}ߏߡ߳��� T�������1�C��� g�y��������b� ��	��-�?�Q���u� ����������^���@);M_6�a��6������������, ��7[mT �x�����/ !//E/,/i/{/b/�/ �/�/�/�/�/�/?? A?S?2�w?�?�?�?�? �?���?OO+O=OOO aO�?�O�O�O�O�O�O nO__'_9_K_]_�O �_�_�_�_�_�_�_|_ o#o5oGoYoko�_�o �o�o�o�o�oxo 1CUgy�� ������-�?� Q�c�u��������Ϗ �����)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� ��h?��ǯٯ���� �3�E�W�i�{����� .�ÿտ����Ϭ� A�S�e�wωϛ�*Ͽ� ��������+ߺ�O� a�s߅ߗߩ�8����� ����'��K�]�o� �����F������� �#�5���Y�k�}��� ����B������� 1C��gy��� �P��	-? �cu�����ڦ���������/-�@/R/,&,>?�/6?�/�/ �/�/�/?�/%?7?? [?B??�?x?�?�?�? �?�?O�?3OOWOiO PO�OtO�O�O���O�O __/_A_Pe_w_�_ �_�_�_�_`_�_oo +o=oOo�_so�o�o�o �o�o\o�o'9 K]�o����� �j��#�5�G�Y� �}�������ŏ׏� x���1�C�U�g��� ��������ӟ�t�	� �-�?�Q�c�u���� ����ϯ�󯂯�)� ;�M�_�q� ������� ˿ݿ���O%�7�I� [�m�φ��ϵ����� ����ߞ�3�E�W�i� {ߍ�߱��������� ��/�A�S�e�w�� ��*���������� ��=�O�a�s�����&� ��������'�� K]o���4� ���#�GY k}���B�� �//1/�U/g/y/ �/�/�/>/�/�/�/	?�?-???�A;�>����j?|? �=f?�?�?�6,�O�? �OO�?;OMO4OqOXO �O�O�O�O�O�O_�O %__I_[_B__f_�_ �_�_�_�_�_�_!o3o �Woio{o�o�o�o�/ �o�o�o/A�o ew����N� ���+�=��a�s� ��������͏\��� �'�9�K�ڏo����� ����ɟX�����#� 5�G�Y��}������� ůׯf�����1�C� U��y���������ӿ �t�	��-�?�Q�c� �ϙϫϽ�����p� ��)�;�M�_�q�Ho �ߧ߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{�
������� ��������/AS ew����� ��+=Oas ��&����/ /�9/K/]/o/�/�/ "/�/�/�/�/�/?#? �/G?Y?k?}?�?�?0? �?�?�?�?OO�?CO�UOgOyO�O�O�O����K�������O�O�M�O _2_V,oc_o�_n_�_�_ �_�_�_oo�_;o"o _oqoXo�o|o�o�o�o �o�o�o7I0m T�������� �!�0OE�W�i�{��� ����@�Տ����� /���S�e�w������� <�џ�����+�=� ̟a�s���������J� ߯���'�9�ȯ]� o���������ɿX�� ���#�5�G�ֿk�}� �ϡϳ���T������ �1�C�U���yߋߝ� ������b���	��-� ?�Q���u����� ������)�;�M� _�f������������ ��~�%7I[m ��������z !3EWi{
 �������/ //A/S/e/w//�/�/ �/�/�/�/?�/+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�O�O"O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o�o��!k������Jo\onmFo�o�o|f,��o��o �o-Q8u� n������� )�;�"�_�F���j��� ����ݏď����7� I�[�m�����_��ǟ ٟ����!���E�W� i�{�����.�ïկ� ������A�S�e�w� ������<�ѿ���� �+Ϻ�O�a�sυϗ� ��8���������'� 9���]�o߁ߓߥ߷� F��������#�5��� Y�k�}������T� ������1�C���g� y���������P����� 	-?Q(�u� ������� );M_���� ���l//%/7/ I/[/�/�/�/�/�/ �/�/z/?!?3?E?W? i?�/�?�?�?�?�?�? v?OO/OAOSOeOwO O�O�O�O�O�O�O�O _+_=_O_a_s__�_ �_�_�_�_�_o�_'o 9oKo]ooo�oo�o�o �o�o�o�o�o#5G�Yk}��$UI�_INUSER � ����q��  ���_MENHI�ST 1D�u�  ( ��p��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1�B�T��f�x��)	��63A1/�ŏ׏��� �~��,95,18���J�\�n����!�,148,2��Ο���&��'����7��N��`�r���r/���e�dit'�LAB_WELD_=�گ��������4ʯX�j�|���p�����ȿڿ����q������ A�S�e�wωϛϞ��� �������ߨ�=�O� a�s߅ߗ�&�8����� ����'��K�]�o� ����4��������� �#�����Y�k�}��� ����B������� 1�.�gy��� �����	-? �cu����� ^�//)/;/M/� q/�/�/�/�/�/Z/�/ ??%?7?I?[?�/? �?�?�?�?�?h?�?O !O3OEOWOBT�O�O �O�O�O�O�?__/_ A_S_e_�O�_�_�_�_ �_�_�_�_o+o=oOo aosoo�o�o�o�o�o �o�o'9K]o ������� �#�5�G�Y�k�}�hO zO��ŏ׏����� 1�C�U�g�y����,� ��ӟ���	����?� Q�c�u�����(���ϯ ��������M�_� q�������6�˿ݿ� ��%ϴ�I�[�m����ϣώ���$UI�_PANEDAT�A 1F������  	��}  frh�/gui��dev�0.stm ?_�width=0&�_height=�10	���ice=�TP&_line�s=15&_columns=4	��font=24&�_page=wh�ole���ϑ�) � rimX߁�   ���ߪ߼�������Y� �(��L�3�p��i� ��������� ���$��6��Z���� ��  z� �6�ߗ��������� ��D���9K]o ��������� #
G.k}d�������n� &��6;/M/_/q/�/ �/��/,�/�/?? %?7?�/[?m?T?�?x? �?�?�?�?�?O�?3O EO,OiOPO�O�O/$/ �O�O�O__/_�OS_ �/w_�_�_�_�_�_�_ J_o�_+ooOoaoHo �olo�o�o�o�o�o �o9�O�Oo�� �����r_#� 5�G�Y�k�}������ ŏ׏������1�� U�<�y���r�����ӟ FX��-�?�Q�c� u�ȟ�����ϯ�� ��~�;�M�4�q�X� ������˿���ֿ� %��I�0�m���� �����������b�3� ��W�i�{ߍߟ߱��� *��������/�A�(� e�L�������� ������Ϟ�O�a�s� ������������R� '9K]���h ������� 5YkR�v�&�8�}���/!/3/E/W/)�|/��k/ �/�/�/�/�/?i/&? ?J?1?C?�?g?�?�? �?�?�?�?�?"O4OO�XO��B�<��$UI�_POSTYPE�  B�� 	 dO�O�B�QUICKMEN  �K�O�O�@�RESTORE �1GB� � �KO��5_BS0_��m`_�_�_ �_�_�_t_�_oo+o =o�_aoso�o�o�oT_ �o�o�oLo'9K ] ������ ~��#�5�G��oT� f�x����ŏ׏��� ���1�C�U�g�
��� ������ӟ~����� v�(�Q�c�u�����<� ��ϯ�����)�;� M�_�q��~������ ݿ���%�ȿI�[� m�ϑϣ�F�������x����GSCRE�@�?�Mu1�sc*Pu2J�3�J�4J�5J�6J�7rJ�8J�'�TAT�M�� �CB��JUS#ER,�1�C�T+�L�SksT���4��5�ԕ6��7��8�ъ@N�DO_CFG aH�K���@PD������No�ne�B��_INF�O 1IB�q��@0%ߌ���z�� ���������'�
�K� .�o���d�����������L^�OFFSET' L�Iu����� #P��,>Pb�� ����� (UL^���� ��O��/
/:/���UFRAME � ��.�[�RTOL_ABRT^/�Y�v"ENB/p(G�RP 1MY�A?Cz  A��#�! 3��/�/�/	??-???�Q;r&�@U�(3�+MSK  �%q�+mN[!%i��%�<�?�%_EVN~ �4�-��6�2N

� h3�UEV�~ !td:\e�vent_use3r\�?B@C7GO/���F|L:ASP@A�EGspotwel=dwM!C6�O}O�O*P�4!�?VO_I_ �G�1_8_&_|_�_\_ n_�_�_o�_�_�_So �_wo"o4ojo�o�o�o �o�o�o+O�o �0��fx������zFWRK 32O��&!8�y��� g�������� ӏ�.�	�R�d�?��� ��u���П�������*�<��M�r����$�VARS_CON�FI"�P
 FPv�����CMR�";2V
�9���	4ೠ��1: �SC130EF2� *���ę����x�0�5��3�?U�a0@a0pU0ȅ�' )/h�r��Ȁ����ҿ��Ϳ��k�O5A���7ϲ� B���R� ��V�޿wϾ���jϿ� ����������=ߔ� �s�^�pߩ�\����߾��IA_WOQ�yWi��v,		��F�(�6�G�P ��I��H��RTWIN�URL ?&I���ߎ������������SIONTwMOUO � ��BXS۳�S�۵@�! F�R:\�\DAT�A�O  �� wMCA�LOGN�   UD1A��EXr���' ?B@ ������`����������x �� n6  ������6��?  =���M��J ��g�TRAI�N��\�Bd�ApMQ����ңY&K (�ѝ	���� �%[Im���������_�GE)�Z&K�`
��
� 
�?"'���RE,�[�)����L�EX $\���1-�e��VMPHASOE  &E�N����RTD_FIL�TER 2]&K �1��_� ??$? 6?H?Z?l?~?�?�?� �/�?�?�?OO*O<O�NO`OrO��SHIF�TMENU 1^^�
 <��%���O����O�O_�O �OC__,_y_P_b_�_ �_�_�_�_�_�_-oo�	LIVE/S�NA��%vsf�liv�.?o�>� SETU��bbmenuxo}oo�o��o#�E)�_k�HM�O)�`.�z��Z�Dta\/
�<���P�$WAITDINEND��!r>vvOK  ꩑|���S��yTIM.����|G}� �0�������xRELE�!@�vvsx��xq_ACTU`�?��x_J� b���%�o@����R�DIS����vpV�_AXSR|�2c�Yyw�D(|�Ӡ_IRg  �&t� 7
 ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ�p�ϬϾ�NXVRy!�d7~�$ZAB�C�1eY{ ,�� ��2����Oq��V?SPT f7}�r.{�
�j�o����j�ߣ�B�DCSC�H{ g�d���IPRrhY�6�H��Z�l���MPCF_/G 1i��05�,��q�MP�j�6 p5������<�0  ?O���{����y4�P?�  3��L?+�ﴊT"�C��7���$����?�� �{����ڴ�|��� �'}&&�*�3\�L2�Q>:����.��F�_����5N����1��h�
��3��������/�� ���vL�KzrC�3���B���B�3�Fu�N bR ��\V/B��^ �>
3� �������,�>�P�0V�h��Ą�{ �k�W_CYLI�ND�!l�� ���� ,(  * ���Ӧ��/�  =/O/a.��/ ��/�/�/�/!/?? &?i/J?�/�/�?g?�?��?�/�?�?O��2md� ġ�7OGL j�pO[O�O��'O�Oڹז�AA�wSPHERE 2n��>?_�?_P_7_t_ �?�O�_�_8?�__e_ o�_:o!o�_po�o�_ �_�o+o�o�o�oYo�6HZ��ZZކ �ʆ