��   g�A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG���DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPCp��8 . 4� �H{ADDRT�YP�H NGT1H����z +�LSq D $ROBOTIG ��PEER�� MwASK�MRU~;OMGDEV���PINFO� � $$$T�I ��RC�M+T A�$( /�QSIZ�!S� TATU�S_%$MAIL�SERV $P�LAN� <$L�IN<$CLU���<$TO�P7$CC�&FR�&Y�JEC|!Z%EN�B � ALAR:!B�TP,�#,�V8 S��$VA5R�)M�ON�&����&APPL�&PAp� �%��'POR��Y#_�!�"ALER�T�&i2URL �}Z3ATTAC���0ERR_THROU3US�9H!�8�� CH- c%�4MA�X?WS_|1���1MOD��1I��  �1o (�1PoWD  � LA��0�ND�1TRYFDELA-C�0G'AERSI��1Q'�ROBICLK_HM8 0Q'� XML+ 3_SGFRMU3T� f!OUU3 G_�-COP1�F33�AQ'qC[2�%�B_AU�� 9 R�!UPD�b&PCOU{!�CF�O 2 
$�V*W�@c%ACC�_HYQSNA�UM�MY1oW2"$DM�*  $DsIS����SM	 l5�o!�"!%Q7�IZP�%� ��VR�0�UP� _D;LVSPAR�� SSN,#
3 �_��R!_WI�CTZ�_INDE�3^`O�FF� ~URmiD��)c�   �t Z!`MON��cD��bHOUU#E%A�f�a�f�a�f�LOCA� #$�NS0H_HE����@I�/  d�8`ARPH&�_IPF�W_* O�F``QFAsD90��VHO_� 5R42PySWq?�TEL�G P����90WORAXQEF� LV�[R2��ICE��p$ �$�cs  �����q��
��
�p�PS��A�w  ��	�Iz0AL`��' �
����F����!�p�i���$� 2Q� �P��������� Q�b��!�q����$� _FLTR  ��\� �����B�����$Q�2���7rSH`D 1�Q� P㏙�f� ��ş��韬��П1� ��=��f���N���r� ӯ�������ޯ�Q� �u�8���\������� 󿶿�ڿ;���_�"� XϕτϹ�|��Ϡ�� �����6�[���B� ��f��ߊ��߮���!� ��E��i�,��P�b� ���������/��� (�e�T���L�����z �_LUA1�x!1.��0��p����1��p�255.�0��r��n���2 ����d %7I[3e��� ����[4���T'9[5U���{���[6���D ��//)/s��Qȁ�MA¸MA��H������ Q� ��u.< �/?&?�/J?\?n?A?�?�?m�P�?�?�?�? �?O.O@OROOvO�O�Ou.kOl�q��O�L�
ZDT StatusZO�O5_G_�Y_n�}iRCo�nnect: i�rc{T//alert^�_�_�_�_mW #_oo,o>oPobot�e^�P~2g���go �o�o�o�o�o�o	�-?Qcul�$$�c962b37a�-1ac0-eb�2a-f1c7-�8c6eb57836fe  (�_��_���"�p�1!W��(��"S��J�E�� X��C� ��,$ ���W���ˏ��� ֏��%��I�0�m�� f�����ǟ�������h!��u�R����n� DM_�!�����SMTP_CT�RL 	����%����DF���ۯt�@ʯ��'��Lz�N�B�!
j��y�q�u����Ԙ��#L��USTOM dj������  ����$TCPIPd��j��H�%�"�EL������!���H!�T�b<�n�r�j3_tpd7� ���i�!KCL�G�L�i���5�!C�RT�ϔ����"u�?!CONS��M��[�ib_smo	n����