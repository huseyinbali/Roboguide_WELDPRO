��   �A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����WVSCHD�_T   H �$FREQUE�NCY  $�AMPLITUD�E@DWELL_�RIGHTNLE�F]L_ANGL�M&EXT- �8 $ELEV�ATION@ZI�MUTH@CEN�TERX SMRA�DIUS@ER��$$CLASS ? ���������� VERS���  ���IRTU�AL��' 2 ��� 
 ?�  @;=��=�BB�  :L ^p������\�  2)�� 1/C/U/g/y/�/�/��NG  �	4�/ �/�!