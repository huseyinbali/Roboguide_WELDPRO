��   ��A��*SYST�EM*��V9.1�0214 8/�21/2020 A 
  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R��&�J_  4 �$(F3IDX���_ICIfM_IX_BG-y�
_NAMc M3ODc_USd��IFY_TI� ��MKR-  $LINc �  "_SI�Zc�� �. �X $USE_FLC 3!�:&iF*SIMA7#QC#zQBn'SCAN�[AX�+IN�*I���_COUNrRO�( ��!_TMR_cVA�g#h >�ia �'` ��p��1�+WAR�K$�H�!�#N33CH�PE�$O��!PR�'Ioq6��OoATH- �P $ENABL+�0BT�f�$$CLAS�S  �����1��5��5�0VE�RS��7�  �AIRTU� �?@'/ 0E_5�������@kF1@�1pE��%�1�O���O�O�����AEI2LK �O+_=_O_a_s_ �_�_�_�_�_�_�_o�o'o9o�O)W?<HW@ ��zj��0�o�o�i�� � �2LI  4%Ho�o��mA}A�o +
Oa@��v���@�A���� (���^�=�1@�c$"P+ �k�K@����pA��XmA0A@�N �����0�B�T�f� x�����������pF}A Ձ}A����*�<�N� `�r���������̯ޯ��4hL��C� 2�lՏ;�M�_� q���������˿ݿ� ��Ԝ-�F�X�j�|� �Ϡϲ���������� �)�B�T�f�xߊߜ� ������������,� 7�P�b�t����� ��������(�3�E� ^�p������������� �� $6A�Zl ~�������  2DOhz� ������
// ./@/K]v/�/�/�/ �/�/�/�/??*?<? N?Qh�4�0���?�p