��   ^��A��*SYST�EM*��V9.1�0214 8/�21/2020 A %  �����(�AMON_�DO_T   �$PORT�_TYPE  �@NUMJ/S�GNL7 L�$MIN_RA�NGI$MAX6rNOo ALxp �V�~ �COUN}TJ
�AWE0�8 � $A�W0ENBJ $��G1LY_TI�V$WRN_A;LM�STP�
��E�C�.�W�TC�
J�AFT�_CHGxAVRG_INT��{�SAVE�YP~1ER_REG��T$WA� SIG6� OP��_VOLTS�����AMP�&A�E �#E_VL � &D'>% I*f$� �_ANL�  p 
$US0 S_CMD � �PRIORITY��"UPPER� �$LOW�$�#$�FDBK�"�RA�v �!SQ_AVG��#�#SD_� CE� � |!E�% �܌ � LIN�!$�ARC_ENAB�L�!� 0DETE�C�!< ELD_S�P�$PD_UNI8��!92DIS�"��ID IM�#���  v1WFt2V�TC�CF�" �� $PS_M�ANUF ޝ2ODEL�5PR�OCESN0�0WF;EEW0ESC�2�2_FI#1�1�1�7T �_AO�"�2I�6D�7DC1�6L �"{2; � CNV� 7�   $EQ��zxODOU��2?@TBd � $?C 2� kEDD  o , � MM�!$D� ��!2 $F� ��B���2NV7	�JBSEL10_NO>JDATA_s@�@� �2WPpG
�{M
�FWP7 �L@�L
 �W�IR_CLP4� L@ASBU8  H $4���R�4�YPR�EF� �U|"ECU��  JB~ �S   $BP�EEPf#}!SCH>7 � �!���`�1e#dPK�*jFREQ.gULSwbSP�0fg2�y�!hyb*g�F�"AI6 �ZCoVG }�hp dD�e�e�`�	��a��dBVB�aZ�EROy}uSLYO]R�`NT�!P�c�O	U\93�L FORMA0NAra�0J3W	� D�cQW�UXWSCCC �@P8JU\�u�sE�IOEX7d� �A�Wfxcc�pS_91INp�� :1�UJ�� FAU�G"t0LO�0I�PD�!_�G]��R��A�p���STIC�@J�R�OBOT�ADY�H�ERRO�SE�d��`S�g�STA3RTE��!TR�0F~��CHDOG_�@�t��0_ACTIVtW��IH�TOR `OCOLL@�ӃC�0�1Q�2H��qE�2� nQ:2TA�B�0 =�f5)$g1��RE��@92�I� �1R��r�%;E7��S�!S�UC*�N3FAILf��DSt@��LT��sABXP��NRDh2N3Px��RS�0�Y� N3�Q#�+3����)D�)D�)D���S�T�`3�3�3NO� ��B���Y�̤�0���R[2����� 91G�.�*�.��<�^� ;���-���.�S?�0��0PA� h������/HOUR_P��o � ��SE�0 �T<�:1HEpP6��GA�HPZ5�Y7�QLENGTH�"� `�P�#�����S�
BETO)F�0#SɦDn�w�x�.�UNy���91���2}!L�8  � �0���B���@������BISPp0E�RIC@�A)$F�SB� ��CURR �Bm4�!�dbg.���������0
`U!R�E}pd0W0������ NEW��2�PPIP�1_P9Oa�EK_Ӏ_R>��E_DBG`���Tp���3��4��5�R��OTF7 � $��P�$�x0*�nfpNCi?� cJ�f?�*dJ�*g?� 7fJ�7i?�FdJ�Fg��Td��TfUP��9�wPCR7�� ��ل� L�Hr ��%� 4��00��2�X�0�À3KIPTH�E�RJ�ـ�K�Ef��0���W	V�2��Eð;0�0���PHK-1��@�� R�M��CH�SPT9L�0�$Hz��SW��BB��O;NLC�$B�2pf4bgF"WF�1t���q�zE"�!� _W;6�AND1o��!�ND2v3vaSм �A� ��M�� | $�0�@g� e�*f�7b�Ff��TfADAP!�LG�CSENSY�r ���EVP�!� 4?p�Oֱo3�$F� r�r7crFa�Ta rm�'��&{�&�!4�&5�&6�"��f��ʿܼ����B� �6B�6��46��65đ�͒0�7w������P0e@�V���TI���(�)�A3T��TX1�'�EP>��\G5P�0S�$��\�O OVӀI�"[�A�M!ܒK5M� AFܥ�^1BEF֦LN d]�����%��� mq `�ePPW)��:�3�6i r�TRKx�:�1�9MANU���qZ2m�D@D��OS�R�EA � 	 �y�&�`�� Ր�7y��q1^0Y6>H^1MIDU��If�!����`�+�3DEQ�w�CD0�!�j=RG�P 4 ^'�ql&�S�������p!&P� $ $ELAE�caQ�q5Ԇt	�E
����<;�r:�{:�0�TVPK�P� UU �uR�:�MU�eY�U���T� ���S��S6XS��R���W�����FW8�dBd��LAR�*�e*�)eO$�`�O$p�O$��ЁQ_`7�gUSh���EC��L����PW{���_O g�#�e �f�eu�)f��bw|�t���DAI$񲄵@Ew~pLEw@|SIZ5RVu�D��BOAR�Ch� ��� `��ap��r{a��r�Q�U$VE�NDր���EVIIC1xD D�#~�JւV}�IN��t�1��q;�MA0�CwpF�IB�URf�f�,E p $,B/�,B/2���F,�O��,BC���Ǳ��TO�ԩ�_�R.@M����މ;RU=P�� 4 Аo�@-����p�?!L쀸�!�PURA�P�REFLOW�OSTi�Rwp�+���A�0������&��S�_DlqdMఽ�Tм�d'���MF ST /@���n��tM�A�Ԡ�f��ر�$����qAD9JD��#NEXc���4���T_P�!h��1�M�b�#( ��8�S_0!���$�HO�!��,�PFL� GAP �2I� ����BJ3WT`�CY�p��x���[�!�y�.s �!r�@�-TOT �@�U�!U�IApT�GWAR~0V���Ahz���r�Y^v��<�KG@?r��0�k��"XsNp�  ;QSCF�l�"( ��O���#^��cQc�?!*�W�GLOBЯ"����� NOT�!$b��IC9!�!AV��Y�\�$"�5�1pž�W_SHF[W$1X#Ɛ"I-�\� ?�t�RY�3`���p�3P�L@M�t���E�NF UIFo�0�O|�p��!AD��\�A�PCOUP����#� @��(�-�
 �5�x�EQ{��@M�MY��T���T���<
P�0USTOz��  ��{P}��w 
�EMG� n�A% ,QMG��,� ��NOѠR�֨��7�����& !����э����s �Z2T�IR2T�qR��E�p�X`M���?�MI�T�CTSK�_WAIII��V�G	� S����7���T�_BUF����g�C`�ABNe��`��� ���������D>�=����GcSIN���R�E���1CT��NX���L�p�7���SsAVH��_PD��4I�e�W� LTn����PIP�s�0BG a`��[џ�fџ�qџ�v�P s�SPC�'� ,>#���b��Aҕ���� ���PP@A`z�����i2P��>�cHE�@i�?! k!k�r��bk�" j���"`�B��� SpB�R�B������_FIL�W�pB�UN�〷�b��F_@��.<�0wp��N�PSVO �C�0a��;PR>DIO�И�`s�p��TMB�^
PAP��� �󞢁_DYNe1i�W�r�F�`KEYe0G0��`@8�BF�1�@���� $#�RPR�O�U,$C"� �B@bCCAL��@`�`T��4i�P�_#!RTy#H���0A����$$�CLASS  /����! � � � � <0S�A�'�  ��!IRTU�0�/� �AWAO���A 4�!� � �!�!;EAɐ 2�(054;52�!?�Q338b51:5J5 J6�?�?�?�?�?�?�?�OO,O;96EXE <
01?C?U?g?y?�O �O�O�O
__._@_R_�d_?OɐS R!> gA�%�_�_�_�_�_o o'o9oKo]ooo�o�o��o��3NLG �2"< �q_qC?�lK<�!A��okK	�; Bд!J X�5� 2�%��c�Gene�ral Purp�ose� MI�G (VoltsK, t�)�p\ ���p
AWMGEN�L.VR�vA*?EGLMG1�x�C1
�rBnu�Pxv�g �q�!�}<�N�`�r����sF�o�hCNV 2�	"<�2����sG 4� ��$����W�6�{��� l���ß�����؟� /��S�e������z� ��ѯ������+�=� �a�sL�=�����C� ܿ�Ϳ�$��H�Z� 9�~ϐ�oϴ��ϝ��� �ϣ� �2��V�h�G� ��k�}��ߡ�����w� ���@�R���v��g� ������������� 	�N�%�;���_�u��� ��������&J \;���gq�� ���F%V |[������ //�B/T/3/x/�/ i/�/�/�/�/�/�/? ,?��J?t?�/�?�? �?�?�?�?OO�?:O LO+OpO�OY?�O�O_O �O�O�O_$__H_'_�9_~_]_�_�_bNV�WP 2&��\�dT 
�_oo0o�d}USTOM 2}&�l  ;oP�o�o�o|	�d�e�nrDEFSVpR&���P<�o�s�Default SchA*w N`������ �+���a�s�J�y�𩏀����RFBKL�OG1 @[mTlaBG�����#��5�;�ۈ2���C�  s���������ۄ�LG_CNT  �[moa�RIOEoX 2[lDEe�A Ec��	�@=i�@=oa�a
Weld Spee�a~�cIPM  � f�x���������ү�|��Eb $?���none=k�#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ��������������R� 2�\
��d6??Ecn���Eeq)������
F0��`^�`�8?���� % ;M_q��������Ee���:[��_��R����� %��/#/5/G/Y/ k/}/�/�/�/�/�/� ��/`?C??g?�/ ���?�?�?�?�?	O O-O?OQOcOuO�O�O |?R?�O"?�O_�O)_ �O�?�?q_�_�_�_�_ �_�_�_oo%o7oIo [o>__�o�O�o�o�o �onoP_b_3EWi {������� �� �oD��ow��� X���0�$���� +�=�O�a�s�������ໟ͟ߟ�@�OTFW 2T�g����:�Տ^�p�G���=���*@�󭯿�~I�PCR 2�Mpe�BH��*B��hh� ���C���!��ffA�  =�R+d��ϩMܠT�C"���R�ؠOܠ]T�#���>��G��C�ǿ��	����2345?678901����AB_L�D_10�>�P�b�B�cϝ��h�f���SRA�MP 2��f�$�����գRGSEL� R� �  	Proc�ess ,�1��2D��7�3����8�4��t�5�����'���7����8�����ܠT�� e�*A|���A@���B�&�h�Ѭ��Voltag��	v�s��<�DywF�X�@]yl���Ѱ�Wir�e feed syp����IPM�� <��M���� �翝� ����*�<�N�`�r� �����������������D�|�' z  �#��E�B�g���o���ݵt���V����ѓC�urrent�Amp�ua��� ?Q-?Qcu �������/ /��h!��h%h!��h!@��h!��h!�h!�, �/qװ��������!��@�!���!���!��L��/8��?���B��Z�� )h/�	K/��?�?�?�?�?
��S3 R&�$��4ᨵ!O3OEM�?�:EO�O �OSOeOwO�O�O�O�O �O;_M___+_�_�_ a_s_�_�_o�_�_�_ Io[oo'o9o�o�o�o �o�o�o!�o�o' i{5G���� ���/����w� ��������я���� �+��9M�k�a�k�}�@��)�ß������a����,9բUPܠ� ୔=�o?׳33:�>7�=L���>;�,�!��"���#��$��f���I�K��?^��>���r� ?J2`�WI_RE 2!�<�������>�3�>�G(=�J*]�SCFG "���v��#g�|�������xO���#�OUPLҠ#���j�,��� ��w>��w;ۿO�������ѿR�I�[̇�NB�  ��� �US�TOM $�
�6c�ɿ �EMGO�FF %�6-�#�LO*�&�ϑ�'A�P�B�M� �uf�x/  ���
,<������ā�f���PC�R ' �e�@�bD�CE�5����� D�_%��M�5p���% ��