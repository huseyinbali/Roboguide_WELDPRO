��   ��A��*SYST�EM*��V9.1�0214 8/�21/2020 A 
  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41�� d =R��&J_�  4 $:(F3IDX���_ICIgMI/X_BG-y
�_NAMc MO�Dc_USd�I�FY_TI� �
�MKR-  $LINc �  "_SIZc8@�� �. �X $USE_FLC 3!�8:&iF*SIMA7#�QC#QBn'SCAmN�AX�+IN�*}I��_COUNr�RO( ��!_TM�R_VA�g#h>�ia �'` �����1�+WA-R�$�H�!�#�N3CH�PEX�$O�!PR�'Iovq6�OoATH-� P $ENGABL+�0�BTc �$$�CLASS  O����1��5��=5�0VERS��7�  �=�AIRTU� �?�@'/ 0E5�������@kF!1@�1pE��%�1�O���O�O����AEI;2LK �O+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9o�O�)W?HW@ ��zj�0�o�o�i��� � 2LI  4%Ho�o��mA}A�o+
Oa@@��v���@�A ����(���^� =�1@�c$"+ �k�K@�����pA��X mA0A@�N����� 0�B�T�f�x������� ����pF}AՁ}A��� �*�<�N�`�r����������̯ޯ�4hL;��C� 2�l Տ;�M�_�q������� ��˿ݿ���Ԝ-� F�X�j�|ώϠϲ��� ��������)�B�T� f�xߊߜ߮������� ����,�7�P�b�t� ������������ �(�3�E�^�p����� ���������� $ 6A�Zl~��� ���� 2D Ohz����� ��
//./@/K] v/�/�/�/�/�/�/�/ ??*?<?N?Qh�4�0 ���?�p